/* encode the mipi frame to send to processor */
module rah_encoder (
    input                                   clk,
    input                                   vid_gen_clk,

    input [TOTAL_APPS-1:0]                  send_data,
    input [TOTAL_APPS-1:0]                  wr_clk,
    input [(TOTAL_APPS*DATA_WIDTH)-1:0]     wr_data,

    output [TOTAL_APPS-1:0]                 wr_fifo_full,
    output [TOTAL_APPS-1:0]                 wr_almost_fifo_full,
    output [TOTAL_APPS-1:0]                 wr_prog_fifo_full,

    output reg                              mipi_rst = 1,
    output                                  mipi_valid,
    output [DATA_WIDTH-1:0]                 mipi_data,
    output                                  hsync_patgen,
    output                                  vsync_patgen
);

`pragma protect begin_protected
`pragma protect version=1
`pragma protect encrypt_agent="ipecrypt"
`pragma protect encrypt_agent_info="IP Encrypter LLC, http://ipencrypter.com, Version: 23.7.0"
`pragma protect author="Vicharak"
`pragma protect author_info="Vicharak Computers Pvt Ltd"

`pragma protect key_keyowner="Efinix Inc."
`pragma protect key_keyname="EFX_K01"
`pragma protect key_method="rsa"
`pragma protect encoding=(enctype="base64", line_length=64, bytes=256)
`pragma protect key_block
THHkDdlCGS49VQPGXLg2qkCU/VhsnuLusCW38DN4OLbSqq6u5iojugI3cTbhvZd2
Wge7snGfPvkzNPUetXxL1J7wAiLZqZrfsRjuJT7XoG0tP8wNrtbC3a9/kDYnopvH
XZffQTdXuLl+3PWU9RRBGPB5paKbRX07SNh11+yh8ik06r6HgU7mu1xUzhJkWQUd
a5qCCBN8zXBdxq0RMoCThJkugIENL6pGl+0ToN9Jja2/N8YEvr7eYbDOyxSm5I55
103jBr1DQUkHl5yHqSD3lyMbRNHAbAvynOlZrYPprLQIzzoiYVj5ES0akwStze31
ZKY/szVyRaD65NvCVEanTQ==

`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-1"
`pragma protect key_method="rsa"
`pragma protect encoding=(enctype="base64", line_length=64, bytes=128)
`pragma protect key_block
oeP8QlO+ibm+yweS8UGA9fSe7tXQaDWu91kQEt5q3ckIDYXz91DEpTyhrTnUzu/S
R81+lUeMX/Q1rK/EDchn71uQdC430UszQBescb3g8p7REcdW+FfAy6w5zEDHcQzL
au95SIe8e8eF9BifEjPoifX7ylStQL1Y1sgppV+M9BU=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype="base64", line_length=64, bytes=9524)
`pragma protect data_block
b5AOb/ftbWP+aUFdTPBaeGO57LwkVo/jkUC42U0oz76rg16euezVXWgQ4wKtXqfa
csmQQ/xj5tszhzdvfP+eo05SUWcsNNX//xgBX8C8juzeaogox0y921r/a/X5dLFM
CeMm8mPW8GdnQIzDsJV4xjVb4evXsdsQC8rqrW0nTFhQ0fzQwsdCKOMsTomqZR2Q
d460sPQOH3AoJKbrNlA4lGyxhRgz5xguIJ3wDh+zMBItsDpW4TcgLhZBWa2u70ST
V/P2IZhrHHSQcP5wQh9COM8zJEk+Rd2QThJpNSaZUSdKu13Nreh+xvHMftGxbq0Q
jZbS4Pf/ZzV9CvVox+HouRoHjpEHs8mGzVMid9bmVnSTi6xRGEZyrXegtUE+3va7
6wc/gSdam50gnpQDbl+ebDZMVjGWBVS2usAbuebma3ZSIn/RkJ15o34/s+r4v1pc
9v7LP95eYS8RRw9vrBrf+9nHe1ohuyF7ycslFZUX6AOSw+OLyog4wmUeWyMZJ0eN
E9knAGL6DD2CmQlru5OI55UoLQ4cw9hUkHSbuOuKIyL/V/dY0u3dD37WKqtbVSEd
XaxRcbMYq34zCk+OqnpmV7Y0MeuV7pVOQpN3YRpQ2Y4Z7PrvIRHKn0bWK3uIADDF
dfgETvwlaV1SJFp1vMYrLke1g9PPBCASwtOrYIERC7OpYK/MJTOm1zOwa66vVIIg
gd+paYm3xhAcuWKrlN225uJvmxYrH++E/GpNrpe5K0mZBpM8088GnZEI1r7fQRAb
iZ7tnDEHUk8cNnOyyQfPernb0+37MCo758yslSIJz3a1wH7i/Er9JDx7Gehm6KVM
YMSvfMOA3N+TuMO25BAnpRnzeYbnGU3m5L3qXuW1mpnhRi+FMM/jutjnoEVWIgGe
fTY75BYUz/cGE5JAdUNazEwIjRst2w5fKvG2Z2L1HoB3GU5Ekpe+U2AYQ/+deSos
rR5+wpo6OKLJXI73zaUdL9k5RitDMSpJIk6NExl+Ri4zEB8/XCYlikRW/7TTtQWe
SKfRteAH4BHnLWAVkQWngPNrJWF9TuWLYy5dk8saDIFrGyDTnWO1LBKl0pE7N1Pg
nM7xSalJmiAah0LH+ujL4UMf0mW0Rq4baddWKUBTHd2j+oxoqPia4z2W1mCzSIuE
Nlwy/WOJPs8GEonzI0Cvw0W4qTLTR9hC42M2XopTO6hHGFTLzHaoHPq4Nufr63+v
d6YDN6Zr2ecOdfZDsRcsisiQcAILlxmiyeoeQWdGRZmv0NugsA1LltEhuDd/358i
ppqrcyNGqVQ4kfAHgbi+dbh4WDFSY+ztUNrDW21SL0hcnBxfCywq4Uwx1p+viBlR
DsjSDYi/7YqFXpSv8k6mGF3OgybByVVOcs3z2zszph3lIr0HBgvkXq08MXwVIxSP
9Ea9G9aaCQavgGP41diT8QglFpbSt2xWjjNgMdRS/5oeTq97C3EkvalgaZHfvXMb
NfIkQr9x3poU7rJnW5jIxCW1xAXysWOzFOzdetTXD+ryXd77ZYaW7cAowHKNNEyz
dVgRPK9E5qEMSw9XRrW8qTbxCTBsk4NS3sr1GdbAi5tXk8A5HRlEVm5dvVL1SjVy
XDjxisOEGmdgfTHSZuzMZ1H3znVghYkLw4QXKVQisRkXowLkkGrJbo2eFoqc0k6d
92fjjKJ82SIvvKVfZIAf47pzW7kEgg5eZYU3/kMdNvNP3pne+rMfwCjv8w1gFUwK
vCRGVKeBSXJAn84EZuM4rLkZ6sC3B2AtP3UYEyolpsUi/wEyDX6UWEMCGvQDVXmR
jeXUJ4PbCihobSFwkrmF3unKO/PdIfnV7FubgWt6WjjLZGcTVzqqxon/eDVNL6sL
MfcRHeoc6opaklGw+LqDo+bfXSW3DoifAxcgQf2nkVqsz/zCI0QfoEhiJ8p9GNOm
yU9sjZYj5VtIw+/OEwRPNM2xzg8aDTf5RE1bVGdubq5DFki+8g+44ti2JMcDMpcu
LQJy/tVney1QDd2HgF/dqpvNsGivfQbFw4r40BWImpmY0/Iz1XoLxhWDNUS6HhoG
N2dOQRd6sctrYKhsgx4UoWkod4jb449WGzPkurQQeE1Gzu4y4NObrjs4B4j7jTMc
sypJ/N1GNebakQoPGCLcBoYaaA3deDuMAwVJLlSK9lk4OL81HdxvQhpDd1KcWcAe
Molxbvn8JhU6rkwP37qNUzZe6Oa8XEi4uI5++RJleoxdTk1XS1W//FTwQ1lDVPA/
W7ry2NqvXIHIypbk98diIHATMqTDqzIF6AwQEBNfYGaCAeHQ6eK/eUshPB9Ba5+J
860bmWvApRwInAO4QxeaJjVEX9Grjjls8ZJhwNK5gP+o1FbBtNLU2Gu1gOEJyEqi
O853etzL9HAFrLq7OvZoKEAY6H5uevX/jz58sbX5EJ3mjJGSsZTox95UTdKzVDrS
IXm5r52DhzqWxBCnSARyb9sVoF7AsUIQTjHfCjRLjq7RNbnNd5Py9fz/UfwV5ccS
/Zl4DGWpJMwdk16EsPDlW/zmoLaJs7ysJYDkxs6oBSHeZQMTyp5iR83XacO+6340
cvq9lhbf+e4oZyar+i/FPZzrZJIriGHahj4gVlvTxQyFQUzVBDfZFIKbdOiN/AST
si5QSvtRjux9q4zYsoY4odKzUYO7ZW6AxxJf+lHf7DWGi8jlzj+wCiec9iAWI8oI
FlxVoMUQb9wp7d+lQiSI9u+qIE5IQlR7t/iJQs7DluM7Z6RsrHEc4BASmP5D7llm
6Qq59jnJee1Mgm0g258xC5xY+w4BnF5i+op1AzrLUqx46Qi77QY5XSpJMU+WeXQ3
RXAFfns9QWHBuPdlhTqZg6sJPYKt2Kxh0zBrT6fkcMzU/CcbyY4zkeBBNfJe+Wef
hQoebaB72tvU6BERebsf1iSXSQPDpy+3eZao4mmHlSqILUxT/VF/tR3eaYuXhCKq
rjQ/auzJg07+q3beBq92h/26frLUxTLcM2NqR6drZEazmzKQw13twjOgf3/hdoBv
cTJBlrwWwdQ6NqGB7ogit985ROqHXNU87sHE9R8c3RdQNNBJYc1EZHyYL2W0fSiq
3krovb279mk1zn1DC9GMPw7V6U0vtwLXejDkPmkb7QJg8STGpaGOWFXk6eKVilFX
d+9e8TuWoThvS1FfPt/VPp6IzG0Fxd0oCk7M2IchOxM2OsmyK4yYMercFt/ZKILC
0DT5AckCCtfPO99e30UD+FAnRskY1/KsH29uRZdhCOuEpgVhH/I9hGyckTOp+SIX
4gdvfh+btzrTBK4Rl8q+vhiUV2hcO0t/bCxnQV3h3A1NruR/f956fd3YJSR7UDuL
nYWxylJEkwoQZ0JszLHPfXW4z9rfp13+wAKDQ8YICANsJb99EhHswOtHqxJ9o9Pf
Ezh4sRcwTEsRllC9M6r74txzw45vrmf0QnBVaiynTYHk/PsCQFnDYPiQgFR3JdMw
XgZgvI6JoFiVTeVaaoShKJUHqLb2moqw+9xsndCUwCX/Em0rQ7uHGMVK8w4hfbU6
nd1pzkw2sKJ9S3PetiFC5LgPOotrOD0xW1tXZRlFSUehaCjGhoI/j4GgcJr/p3C0
Hs5F1rTY52smYHVAwN6SFxhQFXSZTt4Ze7svM8Dgahy1+9Y8lOISCxHZ6En3fDrY
iI9UtvkWrzzuX/K/wmz6NZWT0N2q2TUahfXIzbQdje1kUc00DDUwr0r2v08I1C7N
KlgMwLdckmgI3nypj32L1zw/HGBa7A3QMiHgQSiN0OduJCaoLYY5dm1m1H20G8NT
plge8qor5zxzhgdhJGFb+GPBqtaJ1vabcfcbmOA5r/W3TKdlghbPMToC3jBUfTxy
W48u9Ck+OlIgju2XR5lEfcRmiH7YMdzc8ZQHpo54C+sbn/MYwSatiTZaFdRGn1R2
tQ9ZcXpZ8zPSstUtUa2H4Mg85s81vqYpxs5CXtLVxYRcEVSldK06mi9QEKrRrf89
AQLzs303e1k/PDlfuDuDXpr29fOe2cVY53VySsXaH7ky2OsfL0enrwJbV8Y2s694
NC2Puww6ojhLjNr817AHNCnkEk21dFpijpyF+VggFL/HPpZw4qAwOMToPJHAUhXQ
TCPu0u2HT0VzvJuOHgau/k91Mxt6rEmI2SWYxkr9Yd6svrCP8P7rdYGl7sL4GxMM
Xz2H63KmpyXcQ8QQbTnp7m6rTq8WyX8qEF6PfoTb7gIybdemisj5DoAjjnezTk38
R2rH3aeScgTIssxsxpL1Q307aaYTCqjtIu10JB4OQNXgFsPzXwrZ0Sz361mW89Jw
rMBSBzomh62tlNR6pI1XjbQMFioQtTYYKhUWjs/1Uvj785uMg2xN0QXGB2iST50E
S2DCt9FspILer2hn6DIQpVow87oRWREssAKtv6IBAoVcJIL6YBf43BYHItECBHRb
TJjBElw1ZxfyYqUSvpwRKTaq+sJXDBry2AWH2sa9UK0JssRNddPVI2ORpR/imrpS
uEcWafJMIOYFqoTpoaxjdoQlax4fiOttRDW0a9HT6bRp4dhUA5EFmCpwd+IFp/RH
SPwNEk+vDmXLbsYJKczCHpkVbKpPo8tP7CySX9QbG6GjJ5zUrgmNvwGIgRFjZpbG
vpKj2XTmWjyJMDsW3QWwGvqyJ8OAr5se3XAdwMxtbwpVXuD1SWC4e/hi9J5QNBgb
hZnAcKo7LFt2du/y8KzDDZ1nHe3tgZRbY8ihIUKACF72VWB7/wThv7IfxigEEhBx
CpFlpjgdroyBrhxE7q4b/MyOImLWW+DfHHNeJD5EQ8CHUMIJ5ArAWu1i03A06lTg
Ja61qGIuf7KEbED1SY2ZLUJ9KKNKKODhs3Wye0wYHyjdjJaoxOIGuahaBYFfvoRU
59rvQtz/LzzsUOLf53r6yQwfG9IeG8TMGs1cm1Ph593bgm9V0pD9Pc56W4V/u2od
9e0dXvaCW2s2Ew2S57WfsBmRL4bs1jfFHxSDNGCnxApjALjQjw40a5bdNpcPAdeY
0RnH4h+pqFhbijjTl+5YrEx9zjY/y04xBWkycC/hajAwDQJY3gjfTOyEo0rY60Ue
kCoFW+LMDJr7djRT2J7Z+R+n94imdNtMXOxqx27CzQxkxdqLSWDQ9NZGhID/mCb0
okdSarGPzlQ0KD1ZeG4l2gCw7IMjeb3CKbtGke+SYkxR4J+CRQZa+zN+cH30ix89
3S+QNFnCX3CjQwU+ND9++8F8nhFx5FwsWlwi/FSY5kUv/9h18sXfHzlOKqOxT9cQ
rhILUIAus5zydOAYw9Yst9U/DQglBTuvDpEyARxjIcbesHPd/4oRxgWlXd5HlOG4
a54+rSGyD6A7/YRMWY3sDzdNPkrygqJFfKn5VvujzqMdp+E3KvS6XyaBqVjSpsIe
9mGdg8M2xjsAZ6GM5Xt1QGSBjXw1Ertchx2VYqSJwoJdPDrFx47kFgQtIHutMA0M
hwPQ9X3SL5Gu3BNe3KJ3alr7NxwPmbfoJ/YKouYR5XasImuPgZ5r2qDipm1aEgxo
qlUp8tZnOntvaT14C0bmCcPQxXTztdame1N2gZRKzf8yCzBOlsd24gtHuopeTe7E
5WEEQB2ij9phihVU+ZxRj2Zab/+4k9FeFqM1101o9A4Y/9vxmRfNbivwrMv99HJT
bmq4+8FB4LiqKy9clttK7KqlJDHz+JUpnk9TSvo6YdPO4lXqJ56WMwlhlJuxwiLt
CeB1QuWF7m/9dGstcOzPC9YWhL49ZbkFOEpzZmQUqVOx6VaFH/tKFMmHwg4zl/cp
CvkL5eE1DiAKCcvWKcAD83eCL/dDwy+QWya+w+bxeUFWBkN3NlwIMNFefA6o9NWA
4X3x+UGkKeWWnLB+/tQaPimoRYZ2HWj8CDsFYQ9FudWM7rmotjNl/du+9ZZe4cOk
Ilm9HuR/dttvVQW5paEawYcQNFpiRJWszwa0QSYXdfJf86FhQhbR8al5KFSHV7cT
4N4eGtN7L0LPWYEdojVITei5ZtECDnw+Ew6VtHe/sdfk32CW7DO45e/alXCSjJbW
DhO9Y/UD+l76jkKHHYbILYu/UpVpHgheMO3px7J6lIBmyHAKk5djrr+ds/gTxA+G
oCRG7BMVUUoY1mUVYYM9qIENKZ7HA0EiklC3yCUZP5MCQ6FEvTGhxFox3Nscxo0S
4MWSqZwjGSAHPJqNjoQuUQcOte8T4bSyQ/fQ80BFpCHcCinWF9W1v1Uf/qSi/Wk1
bemYCVz6R+20nnhplJCRCWjcxqsutwYMlN0/xmqLkg8SMCsUHyxywR9+9+pp3MBM
81LmNHorTuY6/T4RLyP1lqjQAUDwePsUdyJ72YxiWrSqo7fmKOzWcGFRgvOz+a4c
NFHG6CRfV4RNkCa9SIlaJR86Xa8/s56slNQsyX8Zr6ih0I12AGovrxhDXpXPLO+M
gbnahs1CavlpBdfVlntDJOUQZhEDReUulFRu8kHF48d6G0HF9eCk8GHvboJhfOWl
WmGxIWu+s7KyDVj6GW9EO4WgDe8GIwhAAKRdf/2qjwEN4lizpbPaRZ2Ndbz05X7q
TaAD+XmQe76MHl1N2uKyI+S2IpuUo1YQ4ToxFmvMGYKeULWqHxzujGbQ+sbol4Jy
fXYpzmgHI5ZdWw8Ie41s7ai5TKV/JnfPD/CSqKIv4RiBGrJ10/sSpzZ0y/0wjGv3
tfE4AgjODzd+OUQxMN4+LFflBLxNGjJrYxkl2YWzRkhSjZMou4lXO7pxMUI5jmRE
rLAFpDkd2JwwuNt8swimSIiG25yBRe59OUuB75AQ8fp79+GlUZfCVqybw3uElQm7
IfH5qF1LcuspDu+qoJjDF+DFTm0z+pcz2pC12kDyprB1UPfzPDMcwyLNDP4RtoRe
Cni/R8bDKlqL2imQvNZXgtzSnKWjdvRj8NGwNTMowdJTYTZpj5mB8RVuYPXrbGts
h9NvQ9w7n7NCtED/SMRfdEmeUULahQLnNVaPYCd8KCSnaIqvAd8fRZYZxPXtb6C2
hjwafiIJVtSjcDxsAtjkKFgEZVru+SguqVx0+XIhot1ozep4ZlWrbpFPRKqNla98
OheaC13ACO5thvznPE82okSoMexxx7zXUNoo0uCNX8ox1sHHY4WjFJdbvOkvPm+P
7J3RFMi5/tz8K7no0dqz7y+zRWdOySi5XB+vQbumaIdPCim1qS89r7jS5jAuW+CR
LtgMkphhu+7+oXERCyW9K+byB7GnfqKLszoPD/lUkCxQ6K8RC0gE8nTE2aHbgPIi
6oS+a+REb5MU3w5QqexzU1TrH/4Owt1N5IG9Sd6sH9pgDMTxd3ZpZ7d5l7GznrRm
/QzylEmWyKURA6Di5QCuMwBfvn5AJK9KSo32Qfm2f2wK6c/gC2b6ZuHMsmBMzdCH
/NyYSf4HMynTiKV6AMLfUY0NNn3c5bwbeYZWhWv2lxD6gqqkdJ/P831nzqZFwDc6
LrBxRYHqjKlLa4rkcHlk+u8PC0deIKaeVbztxNQYecD1d8BE3TSz8A8jt+4B985W
9qrOkVmfYyh7ClvjbMhLRgCnrqMQyXIIXqGJxnSb3k45TPuSIMKGfkvw+dbc2Fo2
qyRLzTfaziGhg/4PQRn+LDdtatKqhdAAIHegbHDbZU3iVGncsknexlplx9LcEjO2
eLg/iVXGTfhb1olCWnyppRRLE80OLT/1A6sAZ41GccYTziroLGWD3AI4rPzuw/9z
aDbHtSL8yULC+P6dA4jsZfxZ3dWhfWMGRNB2vYcOE/p0qO4Q+ZmDNNheyxCdgFP4
5i0bCkfQsgR5tdpf/bomuiW8/7TJvhzgLkG8CMuTdDX7Bw9CgwsDcJvBYp11+a2E
NPXuA4Q2q4bJLhhW3jNkjleHwUbBZVzsAHsTTzyPm+Hy89vXOXbBn7S5JM4GBD2g
NFfTi8HOzfCNzOKKw20zQdecInj6jrmMQ3/AZATVXy1OP9Jch5ZqV4+rsc3KeIjU
bvZZJtALj7Fo/QVtcR7juzoJoaKDR6lL0Vq7d71Zg2x4vyT1SVvfYgdMDWo4a2F/
lMEfnLdtQhjHwUc06dewOTAwDE4454djflygiVw+IdtLqFn1tlW1dFPJyt9fi/Dh
5gPoGXkZGcqfgM2mm7bTjaur5egUKt6kWbu/IjXjOtlHGa+hBvn6CRL78e4WeYe6
afnutxLARwojTCkWH+fJ4RUOZyJY98/jAcJXflVvG3K6/bl0OysdHPwuvDtRZQLk
afX7i+sRIIKtSlm9aviFyqo2WIsW3dXBXo9FaQ5ZO9YirFnrkuL42wwL4OEO8lvr
7Yu2Ua2v/XBShnYe0nVpe9lMIgIxc90xOjdsbErpJLUFFZxkWgfm1YFKlf4Z5ZBr
8qZgi7RArp4t9nwixvaCFn10EBASggagmkq++WIOHrasAV5fMGxilcoJ86onWE3q
g6UE8YmkylQDqyKG5ja/Nhq9z+rDTBITjdclxUCJ5Hfd5OzcG+QwpV840ksBttyB
C1cTpP7jOg0EPhnz30sO4ZZXdxCQh1bcQBc5GTYTbMUpBI6+Gj0Kk1Ad9Fgf/vu2
omJcpVdB/qYn9yi6kPjfy+zKbRpyL8/P0QCeVfyVUTz2mGmnb8P2hwd26dfIgjtA
hmPhfVdbZkSH0c3Sn9AHv7weEb6mV2+02xMkJbUb+sJC+JhEmdtfsMf3oMJGH9MN
+u9gE93goLbZJkjgtSX3kDb7MhHi9nU4KO4WVCLQn0ogu4QHYRfx2TiVnD9Pe169
MQuUEACeP0B3sD1uyAn9PESqQ/9Ij56z9pdGfKlZqun0z2k+xZ1JxaUihqrp7XRB
akmR1S6XdgaAdTY1iUzafbKKbjNyBxkHZihzpzcKfKJYVY/0Kvx0k3F3n1oMeF7r
S9mddQJkSzjIG57JdAMEEyrvZwPBisDbtD1rh9Ktk0HMaLyHoH3xrWcJ/tZoOzBI
eN+1drTUizugw1gL5tmeNFm+uGFVJR8t4+G5swOQ4q73Z5joZQsWj0ZocO/PRWw8
tWrG6rtLxlJPtya0X46Q1HOarMZLFVHJRdvQKCMsXAVQI0FERDc4z+KWtKW49KH+
Rglf1td9B+aJ3EhHyfYypZa1Hc/rQO+xRvoa8cAyfz9Lt88I8JzGkk4otydgu2Z+
gPLINN9sFnJOxRtjdLz1dQTIbS8PuwnzjKQ1Q0hGpfxUyaXVPtlZOll421aUcO75
NqbB31kqwaKUN71uD7aMWPw8eAQ0I9NA4KPQxNeA9XDWfN3rbuwFuBz+NrXLzKG1
AqqBkcqVKO2hLOyV22Ug98anjPBXLIj6Ind7LUozHRJCYp/l3KtOS5ikvqFVfQsE
IitoTTGV9jSWKYZi6Z27RweVA6ltaAVCFJ/Ve5h635DnCcKqy72x0+19XzF4sCkS
gsK873JkB9OhAlLuDeI6rQM9QlYKmsw8jmvCUeP8zdgyNo7n/6q/tlPQnhq8A9+P
JCqVxxBXfzSe2ShwvxAzMLbEuca/99DKGI/O3oyK31VIikZ3VDMr1Ta6SuZLJN9x
1ZRuKWqDhFTz/Y4GowZCxWfiASevE1PNUrw85I6+swE1aW38I81gJQu5CSCx7AGH
cONNgFEXiBZCH1N/6Vgs2YYjlH5bFBeQBiolv38Mn6OySL/Ip/pY5ey4OGAUonSG
w2vWfuTY19FYvqSzGUDeI7j08DL2VXhmqGyemU0B/1UKwHaU88eLphNcBq954LE1
v9j+y3Rkt4hwccn3zVhcbz6oXPHW84PvnVpLmiHY6G0Nu05ND8TA184DefGLE3+L
14NiN0rpX1HAfJO2Z1FXs/fz+O7rwTEupXJpS1KuWsMBFFoQaMqmV2MwBzH1lcAd
W49sbGTQrcq8jXxiCJyrROFfmjfYYO9e+qrI9QMqE3Ld2GoMAI4mZ660XcGjQdra
u8QlU6f6Drt/w93cxdk1LsTOnG0LzWV6/HEEcdzVaOK16Lv56x/K6IpcfKjoxAQX
gXbOW7rfd8Dwyp87UGStlF1RnNsp7mLAYup/u34Ezird7rRXsZkmVj0XxRHBL9OQ
WvOMA7aH46l3xp5H77cze+ugkDsnu9NfT/5K1WfMzqadW1VocKYFG6+TZ7FdJANS
VnZzKaaHtTfGD8kNnsF7W7+kDsTNdiqejvINjR3RCEZOMeKQU3kznI/yv6GFO02S
csK1GjzVzFRRxEG+PtuXhzPAIhY6FwxO9fzNmO5v+A3MThGh+nqLUskUa7740lTl
k8Vly4ls4sEyduRAteN5okffegHCRKRZVz/nMkUgwxaAQAtWtT74MUlgcDeoch1D
smRMa6qIdYHROXjGNDU3GVT2UZMm8YEHEX++Y3rEPMhVSoM6oC2cL+XF3eZUbsFP
781D5dp5BFfgoMLTYxO+44IJV98K9x5q+DpkbxnKWIc0C72dgciSgFnPfKdHcnf8
44PrBcnLVcNLYARkbaYXVBekmws9OsrNBpzXRKBEogrSHRDHXRPUk+c/JezzNFoC
cWGqiOpwlFAxZXr4z75Hhv7W1jcJtHeQpYiZQjt5CmQT4pLxhQLcvBFrdKbJ1iJj
sHuaK5KlGjFijJcuJGDZDdQRuGW3IVSSezwnyOwG0yM41AS0iKW1OOUPbxIvTkHh
5Cu5UWspsG8oeWCl6fzNuKJUxk+IJbOSV83Yr7PzgIgVbmzJk8RAWOi8TxGyYpIW
o/dmzbutTrgXrpqLkVvCpoE4VahK3wITex7lEHZWlXjPN+e4DZ182kYEBeuyPU14
G1mDXmHIKLNX0YdZGUxNgs2XFhXxz0zGLoJLlVjWXlbdxZgLfNhApLO7MiiFMKaP
Z+HFPNAZZM1Bs5FYNdqMuJ4/pdoCTUww5A6azNmix2dHxvafW3oSCS+FfRublN9S
HZl/qv82f9CUpuQfEA0U+tbfw1S2DBsc8+VEdWP/yIFEU6xp/e2GjvllSSmfycms
wN7lDoWcgZtE47OrmD4Pk6kE7L8XscjcT+I25JIVB5MLs8srHmHf/j5fmSznbO51
OEZuH0eZ2hAPEfjGy/f877gNXecT5SIg2124bztrHzj7aQalHNhoghE7U8LE01+f
igXs9tIzqBdzSJUA9QrhpkAuT6Jg6bmZmPC6d561lQsOTAaDuqSrR/bdl/isPYe3
I+9fiImGS74aCngZ2abofmpqWlNqiq6MqBlEpvLZe0UVYTWWETE6LxEV56FnJcVM
VsJ80N1GwwA66KBzdupKM3MZgQPTDIZpQzxKJKswGaIKHAt3lAHI2bHPC0myDHYv
Z+ND5C8hlbE+FQ/z09kXhfcuHQnFu/xBpI11Fv+KEd2Y/Hto86Prb6KG6bCZExVH
GfYjHMztyl5NrPSgRabmKflLxZBP01z2a6QWhh46W6IRYYEb0IRNJs6lvs/qdspa
pBFOZ4ugo4rfVIOQ9qCTLFsvb9i1XqCyfURBfDBBpLP8KSmPjNXGqvnj1sntLxNr
aS22+alVZddmj+9oGoe4DZQgEZ9cxdgIHP+wjqAfFzx3bk9KRBxTZchSAENuZoGd
BcMR4E7a8V4I2Rl+auEwunYcCEhIBR1cvcwE2rS0cB+zO5vb8N5nJHt4ujQbrBmL
WhurQYAhCh7DPwzCpFRbemBXjJtRKsw6bJgX5yxe/kNL/uYJEQgu0vS1r/hRGgG/
uWbWqFDmHIOMkc7DfRRfRQ3eeWhAFhmgU06m/ly6TZvcw5Ap5T2AppKtl1kvl6ZK
keizisMBTP7Pplx7c7ZWj4vbcH79oOMxopVDFt2opiaTnyyUJaOD+tGstCMF7Aeo
+miTOWMWE/YK8k/WBn7QB8iqmZOxxe55iQejb15/1n0WcfoPoRPRQZ91x2WVBw9A
s8uT1M/Zog+anEV1fxvrKEZfwvFNWHzHP64QnwJYsRqJd0APoVOrXpq73LnRr0qp
/VkqeuoTRXbVBLs+8Pn/VBQA4zgjDQnqOyjT8R1B6BymoNSd48mE88EEFev1mYF3
cj4Y5wuCJJaC0UBmNv7E6xBM7hhYCm0bxdcdYaRcLYO0nUjYqwv+qN1MkGdwauxR
00xfW50LSImwZaxogL7y9txtVuYLETCR8NXSuzfb67GPRNnpNSkrHHR6xTG6xspj
KEraaNgHG+HxzT8vLmG9uQgdd9cv+8T0ePzjgCVjU5NcJ8Bj2U5Q306LLxeu9y/x
NCUUcBhbRjk33sa5SjjiOWLL1Yd5T5Npo6gwwoLKZgjdyDh0xrO4bf/glKOxuCnf
+XmXvUGloMpX5gVcKxmmlHP2FZAxPGXuC8Ie87B9j5E3/purJhPhJa1pLXZXQRwP
XQGCBmq5Zzz+NZtAoNSGZHIujiinQUJAEMeYIeYwV67infx9Pzkw0PfpHR4If8ea
uIrHbwxilNfr+xwplt1kkQA5XU7nClD6oQ/VPbMClcO2u3Fwgv8PRt9pK1nvnRU4
ouFoxxIkorO7ornxKhY7LlnzQthzJPIIRElurW+oQRjwVzokdH1SUOQQnvbLxxFf
P0zmdpUWSxnWuLrorRb8+qyliqY4bWFu/sU/XKCRxrVWhWwzUiN3u9zRhzI8f8Ik
7rgNue9Ylx6Hg55/hit42aThcjsBAzLSWcwe+H5+95ua1lGJYgPPV80WJl5kQmNn
TH9oY/7IS3l36hQIFqQJZQ/Axpp8zcjkwd0h8tCR28fU5+OHsMA2PaJibcC/t87X
YwxcFz24xMXgjBWd3bRRtmAWJf+N7V2IswE5s8mbwl+0NUQF5yJO6ZO3pC8KDIWi
kOGxeQ/PyJeO1fat0TL68mTTTYdoeDZs/KiyNnujEd0=
`pragma protect end_protected

endmodule
