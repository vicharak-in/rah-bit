/* encode the mipi frame to send to processor */
module rah_encoder (
    input                                   clk,
    input                                   vid_gen_clk,

    input [TOTAL_APPS-1:0]                  send_data,
    input [TOTAL_APPS-1:0]                  wr_clk,
    input [(TOTAL_APPS*DATA_WIDTH)-1:0]     wr_data,

    output [TOTAL_APPS-1:0]                 wr_fifo_full,
    output [TOTAL_APPS-1:0]                 wr_almost_fifo_full,
    output [TOTAL_APPS-1:0]                 wr_prog_fifo_full,

    output reg                              mipi_rst = 1,
    output                                  mipi_valid,
    output [DATA_WIDTH-1:0]                 mipi_data,
    output                                  hsync_patgen,
    output                                  vsync_patgen
);

`pragma protect begin_protected
`pragma protect version=1
`pragma protect encrypt_agent="ipecrypt"
`pragma protect encrypt_agent_info="IP Encrypter LLC, http://ipencrypter.com, Version: 23.7.0"
`pragma protect author="Vicharak"
`pragma protect author_info="Vicharak Computers Pvt Ltd"

`pragma protect key_keyowner="Efinix Inc."
`pragma protect key_keyname="EFX_K01"
`pragma protect key_method="rsa"
`pragma protect encoding=(enctype="base64", line_length=64, bytes=256)
`pragma protect key_block
YVNrsGvh3EnZLrMpO/BLxAuuueCd4qNixgKwiSOCNHMJU1UE8Oku9ifgQgTIUttI
LCx+7qSrPNF9SbhytB5u9YKeSJ2gRJX9X+plnqHOqeDJ/Jne6kstQ3HPOyr1d8N4
5egdj3Nkc+Zera23vCCUmoo/A9Pn98ELbEn5SYY9p/Ue6bHYawozJ5TlFIignigY
eICpFIIyrYFxdCyJwO+oR/UsuMeEafo+ycUEzNZYL9n315GSo2uvP6ebNQZNUCL4
tT8FdPz10/ItyCTKQszUrwncba0rtGREZYPBU3fnDdys94xWXpN6pgCjRwkosE8w
VhPb5exvrinwiZHk2GvY0A==

`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-1"
`pragma protect key_method="rsa"
`pragma protect encoding=(enctype="base64", line_length=64, bytes=128)
`pragma protect key_block
EZ1ERrzrOJhMfOGbPw62T8WPbZiJxLdrdKifvSuv3+uuySyxQuAoEMeimKuhujnD
TT5990eVw+d/ckpHNDtAs5epbajI+Lyn2zXmqWvNnUW4O/2baRyTY+yO/xE6zMr3
RuCKFWXb/1mUMovaT6OpprFwagJEKNI0PaAcsepZsV4=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype="base64", line_length=64, bytes=9634)
`pragma protect data_block
eIejs49xrXI4La+JRLfgG1VzBwchR6bmcain6+4z4TkqhWvlK1zBvq4LyUBmY03j
ZCXRI9L+5wZu2BqBgOkZTuPIZfEjrCzLb1F8idhEl4anbmTkDCU/cvPzBnW4k+0Y
hd9MlJvaPBJBCovdzLY60Q3iKnsX7xnFSPRDe74xZSo0+22sJVO1o9XsYlUamjCf
1cs7LOcdVJhVUiM9XgJ0SWx0t47uOhb+DcdPq6E2DmMGVExKIAFkNEf7oOK3YY6w
sC8QdzQpI0RrGfVEop9jYEHvgBwmOlTMtogvRfoRBYmwcXHhqv2BWjkG1qv9ZHFq
qU83uMpk0FeQX7wSx0JQTnDo4kR7co3Xy7VG6fdlVO11FdCKq85Tf3p6BM6kD1uu
YzI8VXx2wJgRKimLP4mGgJypMxX/cubTjbrE5ESApQrHTE2JAsabnj4MyvadVbdr
BEgchKr4jHO4RT+TE11KXTAZvsTtMOZ1l1nKlittI0YcuoGrwXED8IgxdjOKMyDl
Ysxu1GGMXxPpmPwhfVI2mocx1Iy6VQlFiADtr38QXIlrdFNGRHXGDva9Wv/MJ/f5
fEiIM9tJMQPrazlrs49F0QAjvMzhITbu72BKGfWYv6KPwr2LZ9jhjFrKoVB3XTwE
j+/0YKNibgvW6nqUQFSLjFMBfLJUmhyFIzLFCFBiNy6KQVx7fvk5p19Ye930WisV
tNrxTKcF2GaU0C1BPrxOI+QtjmITeAjJj2Roj7OmmSpQYRUs76QWN1kDxZv2vBD6
0fMB1Kg5L+PmtAj+c2BHulim9LFARfSEGnUVhRQ7eebvqxQVEXb6n1U2CRbJ6NgA
tG6Znba0E3Xk0wtTwixwdOpqWsoDDCzbZIny7m2kKS4osZW3j2IFvJgPCzb0Lwbw
SI7KzEVee1Mx1Co0doFw5CbhDJizKIpE3onCocrJTlmGZJwmVqbQasUTF4cDN7CF
EfsSmjUg7ZTk4MlZQBN/vaTnhGOHa7zUKhES1CrkmBE45jRZPLgSPkLcE18Iwk/y
jxLAhO+HiHSSohpLk84pvlD7FpPbyykCRKlHBNY8aZv/lofo1BoFxQsQ1Q69JjgA
R2vth/LLf7EQLjOXoSH3ZC2ZqsrhsWIbZH01lwmoKZM2IE+GiY8+ft4kp1PJKl5j
fCKxwseZ8OcNUsQgn8wNri4HuPYEdASL0BHBE0ZnYKdqytSV9Zb2tUQ4D60tvqrn
zpMCVIwpTOlossvtD1W+vRXJDYZz8Q81XOmZEAMaxSLy7k1HL9UXv3RFT2mLT6y4
iMWzZeyQEnZugA96ljRtL9rH7X8VVgsQ9MKBnikcRSBztcAr/UPIY+RWPt1MqOeO
DjkqJmS9+6E8TeI1K4LI1Ab6D9OY/bwEo5pVaPLgMBzMuJJ31KeFLDbhfyBVzPgn
FBlicEIbe/GH5dw/Uz0YIV9SQ2jdzjb5NUW/j1N+A9GDbrudOotacSAVH8BoEJd1
C1bszyARA+JE6HVk47KwKK6lEDa6nVT+4fsgVmliX13VUvjF2kOhd9OnQjkiwEjN
VYourdyDCB6lAvpAT09dk/GWhgpa0a+UIPYj6tTjNMYDk9g4FPWsDlZWXOkLIojI
T7CTL3xk8GvXXA92ZXPd0oEC6za2z+C69wGggNWB5pjwMIi7J9WNGozuF5VX6LmO
jBOu0EOGLJBrfOdUiNEeX3HE0Gtk4lOzttG8SB6urYd2OdOS2kImcd/aAQd0CEaW
jGbT7XxZe4gx8/Q6mjGrI2G+0AUwRVmjPSdPakKMCViyYXPLHx2SAceCBop3+rUy
SYTZYaiTCPhbW3u7unIcRVtHLCSW1J9fC2rrMocZPqrDLtiiQSJFd2tJlXaUgasj
dMMA2wFhBIWNF4UUtHVkJ0lmKG9ote0QfKW79qStqx7ILjSNlhLAq2zpkDf+A4ub
LkB13HhRRTARJgyy9ipGnD0Xfpj+4ihrZOxvCSeGmE1S/YrJAJLlGw+KzpFypuQV
7kJDFpT4KZqUTPrxG8jkRxxLtd3W+U3EVZQywC1dJGFpcjQBK0btQZct2ZFCj3ox
VMqmE5VKzMCfbZyfqIZDahdDL7VfOC5PvJ39/itHQi39gAyRHDwPmVsv41A9LaxA
Cy58UvPnfP+uXLNQTxpjGgWVtAyP3klabOGtqsLUweGghFgJZTWG188x5Up65WDp
Wi6PtbVenWHm5ivNIiv9bsA8Lbe38brbzbKayfZhXHYJhrx3QTN9ZJucFdCBmy5V
zbtEAmTlvRfVi5JXPWADMjayIaK4v/6aFJeeJT9tQ2Uec9erXzRlZwITRfWjtRhy
Thj3d4AYmUeoVAxh6SMXDPducO3EmKraT0osulrBifOKv0Oto2lvnLyDQwYFIgYp
207Em8Ygg/yF/UWflaabi8ii6xA1m3rXZdq+JZkEPtpbGY8QOa+fSkAlloozKTWw
gYU8NxYWz8DK/kwfSnYXT3akVXWIK0nKXEOXvc5B+kqQVbB9f+kZtxNgOOr1VYB5
2cDx6xX3Sbm5L0vEs8LPf12Q1Go5b/hCwhHAr2IYqj7Irmp/Hz8RXY6yZYuleP4I
6f8BKoZOOEI8gEwhkzRBKdtDG042DlGNeYo2q+QirbUOE7VdyvwW0vQdCyZgH+Uj
tg391yHpnwBJKavJ47lNcWVlQaQwYb3JfBwYBUOY1LCZ4RJsnPjQbiGiEkwSx+VS
8205ARcYCffg2MYZH3t5IC1HPqx0OGwks7SORqPxxokcmww2MkXpVLulbMroZxub
+5Jj9ek4mnxBS9Ovd9cfYyLBRGn+lZOMBBC57NAEdWNobWeGj6K7NvimVnB1M9zY
bmGDYLKbicZ5ib1eXZe98r1WuwFPrLu0oqy/KoRPVlW/bSFWTGeLIfwf6Q9/yznX
Ns1lat6OwW22zXXfoqUIdGUeRXFjJbMIC9XUmXZB/1LBtPkXTZhQENwCGG1S3Ft+
eokCtKXncpDZ6HgVEowIHMlfl7utADx8WyCyXd3aKZRSpSyobdSw9E1xzjeMF369
8xDIpxwKal0nDC7QJTRmQTO1+3Z4QFwf0QUfN/KPTUc0vmUixvdKKwCS9NpxFNTv
6xOyONvKhLntUVQBQ+E4w8XClF4CcCSx/5ctdxQowpnbOnVep+dxL3GGJPpco640
fqIuxxrBydePJvs8YVWCQzn9aQ9QcZElwgnmVs5hTJG8LPmF+dLW/y0ErNLenQrq
UjzockwrkTADSFjO7IhZgD4gfyIhCMdOmBCJ6/MSmyAVvmvu+ljcvdRDVYJrl4Y3
AQbce+d4iUhJ9BmTQJ3mFJ6+DibXLh0RlfbAshr6CxNZjrOrHEnRSsiJM7RRVFKB
054vHnzXmLDltm7ZYp5sdKKfkldELodpKIfh4vkou9zBlIsf4gcXTUVloqrBi7pT
u3z977nw0HCl3NPlZrJksIVdn1PFBkRxEYdF/LZFWrLyExqv1bghmdGqRjPD8Uco
u2N1rETBLZs55dMCJ55R2QRZOPpKGxUk7DyhPgvRVR1nXzcDpI7+V7h2XhRoGLT2
K3u0zJNtec3QCdzxWfngaAZQju81sAvVlKMk1jTUJYk6iomzXxFC91/8wPVE9lwn
4iQmX9p+t4G5KTBbEZYzcvxmmhuAQ12gcPQZZj3YQ3hs2A+DnRvwrloOMY/2fitQ
RVhDH/6Yf+Ii2cl4upCrip3SGYKeDry/QoqmEnu8ncp6ATcrEFAUi+mx1ZgO/fe7
Yba+XLufwWBnQ1YCUTsS3w0mAIUlLKkUBYQxV2Hc9WTJ/HilB9Zsgt0Iwj7hSv1L
Qf8tC11ReW3C/lhR2+JVcSuggAxIkBz6kQO6uUCpNoM2V5UXs+G+qBYwwdr8NEpf
qD0dWFWjoHO78d8HtnrWgRK9nO6oEPuw3netGpbI3LP4VdJ1zbQrE6vNnKxDW1WW
5l2ZtWtrOjnbhsxl5/IYiZIUFA/VTE2v3q7bLgIMpSeLvhA/XYp7RgJs9p8Q6g1E
sPZTewOaHy69uxa7SEbyghbaxBCmAnMUmDuRYReDNYBLGEQ6mCKYaRygaKTJBUrr
+eIdu63emc9ou5L0hq9C6WsNaNObnMMPDxHUNkDahq+QJTyAaBpTC0eFZrezR5Wl
cFxT03NvxczqEjcAzjbivGvTQ56Rbs76OKksyhx7S5mEFvyMiuqqtTOwycOK8Zvp
ryfc/CodWY3beHanc+/1KHY7XL0k7FMW4HaGyzm2X2AyV0sC+hrxAe0lURjihYnp
MOOp+AF9WwT6eOjfhm7SOFF9s6FXgQO+jI9OGrG6b062jnk8OsiiNIYJO5WJtInD
i68r3lRccxWwolfE2ztxO14pji5fcXhrUBibgdUF6wXYGtoXh5VTXcIhG2dcue+2
74H2EtkfV02BeiPcSNPkiqyT+r/B0/mRvaqIm6q+GRYDR1qUApbzJCgpzjNbWiuE
ACNXEtc56yNSyCiU6BR5t0hAFerstlVDKKyhBWP4oM9jbzoHb336ltYaH+1tuhHo
1m2O3ZuHoIBHLQGTNBtXnw+tX4QXJ0XI8lkDyymf2YLmvOWiqd6MndX2J/2lTMgP
dEevurVv9hRU5HPmg20jl3Ut2yFhxSp50UeXk5oIbFmd/h91RPiBZaHlbGWopOek
4wwfkKPtoIbrMpb6cFzncuL5E/SfTMA5VdAonrfCj7G8c+rM6aalLOEqJ84+CTcE
LSkxghyiVDX09wF9LuX7Gv4OJe9t2hxLtccjG7U935fNO+tXz1UhRy4Zbo9amurQ
NMD/dvWwRU/BC8D7cGODDouS+J2MYKEf9xKjy7yZvAjHsRWw5gqy6m61nGafWPha
d9GE6FrfH1YrHm/cIloGsrwtQ3Xzr47uUDa5xUMRzB6D15Vbk/eJrt7rlRFWGyM7
cgBBWovlTOChSqOSA9ym6wuZX04ugit87Pn2SMUI/z6MgUrjYY25HiwBYTZphPJm
ue18KIU5KPFxWLGLiGOb6FJpOGwGRq02fB/mecYNV6pWU2UVJx1uWhu1q2ElpFYB
rA01YBduUS8t9P4AnS2/9dQnShlLllbDa971VGyTaqH6edIlhoTh2MvdMWpCBnNl
9LkUD9FgxWGf4tz67zrab47u3mLwyM2mzRAZ1iv0Dp+OhcBDtThG/2bJb++3D6ZG
zefnCXGxFIw9tWosjYoqzOd3aqCR3gIV9m5QLqSeZZ8284rKGXUdMfVRbfBKufGP
d+zfIxiN/42Tj7QBIsS3sXVym3rqPVXK+hZAxofSaPsnSgRp+AKoE3PGd6+ni3y3
bnLWKz9syUA6uCbHHtJgKgL3hDbLBLdfLskI7nHF9c7HrQlKxXX6nwcXT1nflXoj
4JmduDw80QB1I7NUrCw9jgTsjPVKCGRgUekoZS/1Yk1uBEHkZjHBGFJ4tP61whe8
mt8C+/I1w5WKxUveByVHA83VUOGr0AG/T4lQuYtIn6gvGAYpFvnj/iBGDb2KF0vy
KRotKvMPD1OoaSwAjCLaTjd6paACMsE/JjQHapotCKdFF3T0mnRx7tymbtemxz8O
wJbExHleRY0ZZ/oplf/N8mXyMZoZFvUNK7421EzRkzeLX144pHv8rpTV1ETd79U7
p+4oLWOVLithucZUcfoYGXiUJAVGnlA2nFVQXAb038kF7BjqobkeRdcle3dSVtwL
HedZ0hHi22VMVtiW2B8RM8GiFjjceIAtYvn/FCmuE5WltYYk9WCUthBobP+D6Yd9
C66l78ymhQp2GnwQn8cewrkblGW9jWLFw67ZJkWIUv0qWp2+2WgHP4kEGNTwgsua
6KaeEojDQQVIEfrgB/mooCQb6MOGKCg7DqnIdmYpxnd9RS9+3lxP2UfeF++PrxqB
Rky5SSSTvCALmPgSIeKkxfpXsuWeM+gWGannzfTq7fr6IY33NTzQhPsVPPnKtPAK
E0hiebegnzvXhFUww9dnGW9R31XSDYskxVmW4BIGIEfWphV+CDRxW4oolLMT6Gt2
h2SLQ/lBvZrUan8v5evBgs29OPj9y2GtkKJZl8UDjpuKDG24HJ6hr1fJrkHBImd6
ZtLTsf/Sn67nEhpkxu8uwiULBo4SbZjbCNQGor3mJAmEAL8M02wui0tv+P+HuOLV
SxPBJk8msIlv0tPjqqM0SWErY1D90LrGDhhjLe7ZUnzQmam/TF9A2eetx2vEpbKE
j4FS1kB6PR55qyMq+Dh3hZE5DwwXkixibdUxNuK0xQ9E3/cPYPhcwcaZEefPzwla
lJ/oqbktfWoEs5W7g7Lg1DWoEhugamvLyUE9VzvUQFfbveHqNMxfAKM2cuR6zDnV
XQpeW/nhszLCZJ1RLF2i2jJeMPcOQRIFxJozMebXxvgh3Q0VKAaM6zGZ4zDBQpsc
khLV6NB6byo4JturJIW/KEvZCXB5SjQ5J06qF+spXouEFzPNpO8PSIwpcI8jXBhF
/3GqlV34GnwMPRNhZPUpatccOhV3OzUHhLGH13uBKIjzLHXyPDgMXEppPwgT/Zmi
rb1A9Ev+zSQObYGSlQ6cwQN+uVMN0qOVyBRgztXZ/Lxpg6ZG4w4on+giZkScIn98
kWxto12mMWjG0ZT3H6wxTX0joFnxBpHvixIQyp60zQas3egucTvL4n7J2KZbepKh
5QYfeZ/sTCrWJzhMGpVcV+YOYNnd5by8i160zajoy8PlcylPAeymNJ/RI5sPoW/7
hJd2CqmCaCfQ9rFYEugwZKBSQqp6nOqyq86qW30BkeDOqBg3W3t9sV4beAS0jYcI
Dy0E52p2H+FijwAipUI+lR2iv7AXcYoBnkpEzBdnUSvgmDJkoNCeTXDYGNT4IHYc
4N2gofs6GXGyX39YQ2GSK86uDuYAY/ew9934F4/5K4bQczYAS8Q+eZyi1iYwAPa1
rfB5XWxC8QGhaq09mF/JxeHbfhE1Ge38+Qwzb4YNEypVVGcgUGXc6eimhDGThU3d
HJv5pQkbZ7a40gEFuR+5D9eJwOONoK09bOgMeoiPr1HppLjoe1INLzUhj66kKR4G
TyrgqvmY82FAf5wLkUhf8NBGvcYE2S6a6nnX84zbt3LFZs/irrWA92Jvs9Jo8FLo
3HEk4j+8HsYohkfYlFhBSC6JY2X6oMEAzwp7lWBBgEL0xhEokwXC2uFr8qzMwUWo
2qnacfSLv7dZyrR0gfBwZSogywloEIp4UJVUulcDUJnPx9Ttpj+Iye+Umal3UQiE
xhXUXfcplhaUn0LEjl0NmUJB6WwZDHG0UYYOyGxTnn3A8VqtqhL+nriLZW9w5CRZ
Yp2M1ABz71ckyDpTSEu7OERiNbWGCzWOdZZ/6tsGHJqid7G0lCfxLw4gWiV4rVBz
RCasppEqgwrilwt6iwgBQA/VUyn5cC9tQQtK0pkUw05ZCOqVoKX7rikYLLU6omzR
momTTPe5q8pchdjZRUvIA0voYzRuMhnRPhZ7eAWI8jYabUGPd9YzPbFECDmVf3j7
tlOBIyy5MmfR2YY+wZt7jabrR5eDjb2WcEm2nvrCm8dZQU+fMq7L4p2ojKhaLhoy
yHXiBNJaIT90bYq2ZKFvO51vvv0G+9JvhSQs09I9hAZS7PHEss/HZER9kDE58Y9v
kI9UJjXGK9K4A5/PCmGl51wa6r0DX830oZ2qfDpynZo8v7srM1Q+c4xsTTRDzFR0
8HJwIu9G8t3vrDVlLkuCC7iKU0Mx7Fz0l9cv5jK08XQSOa0ZaHgQtWrQslKJBZ76
h4QSYL2+HUPiCq7dvrAjMS8lxMqj/gvirv0hRFNjZfaCNbuE5TPHVt0UXpYEmwKS
45G0kzeHvs3bMCWWkpt5EqzltzG9LJpustHqsV589L6iUs8v5waqw5CYeH9B42zy
B+biZO4rn+RnzJAZTYBFkH7KBj+vpozfBH9ig3WWirYnDY3uRJLQkpHzEAODJQ8q
m+utwSWbVHX6xmw9RC6ydB6RcPIKFUUcTVbQyP/6zAjVg5jwjNueqnxqMhVoGzZu
Om2bjAwPNjayn3EUu7SSs1ULkP9J2fBMrNmviEwzNikwq3OSwQRnG10/Eqg6baYw
LG4R7B5luXzbRkefsCuAgh/JVjiVamAlYsztZYmMw8enfGxNKTJGuqe5f9D4dAD1
y5wASdRxWgk2q3s1YqkXrg5o+OclOPF9I+9Vv6qlFdJDuD8QZ+FUCOAPffEZNMgG
lhZManBx5EcfRVbhT/VLKG4iU4LzQqG5Hh61B9IudIlI+xSRGn+fKxPIu998Be1T
h8M0DRRzsBQl6slxC6OBu85G1BuLaBlIk3z0GZxwjnSftYiJDHIbOrDmXLvu/vnt
YQb/IvxhFOPTb6vpZh/ph4AL2X7XR5PZOdeWXIu++1WT3kH5k9ec7siFtP+wWZFJ
RWqftVcTR7PnROKpjSwHO2OruSUgb1c4QsYjOvACnDg6naQOJRwIKFIiY+XY1rYk
blGmxhY0gmMMHY5AWXAdxgBQiYDzQXzq93giKTn6xYeBDXdgjf50R88jMLf871zZ
+byhjS4w3TBj7F/M/1MjW7uEebfDuiYabtCvunHqANklTC4sj0gh9sh7Buo9Nzls
WR86Fd1rgDrZI0UpIBliqrl8ii55c8h+3r05C4Nz/j1tiHbJyPw6Dg6h8EuIR8lG
NFdNbtzpGZ0sBdWFc7mjnOoAI3oTdyt2T6ix3p377NyWH2de1W2k+D+DAVsofVP5
/clQb5iQ8HGCivoYOhxXwi0eadwlsXJnR1EcSzj9Swp75uxfte0N6ma1NX1bsjQM
th2FiwJRNpQcUkAT6J1wBFacEq3Nu6fLzquw8AOhwmXZLv5yeVZRaDxUOFzyR7gZ
JHi5MYLiCoW+LnDWZucSqRxletFCddkhhhVaPtUJAkemh/48QiSfEaZU7FYjZydk
cD3qgR2IgYxctC3wx6R/WOl19khqloJw1fNeGeuMgiyY/vnAhrvXuinLnJJ+Kn9M
I9MkRuVsuQD+MFp0VXhH84/j5dcMB7WoxpJbvmVx6YvC9FuMfHl7dzDibzWuSLLI
D08G8hR6Hi+sBwIzyOIcmvzaAwh/frue029o1UdXQpe9u4Baf2Z3/PdayoicywBD
0BrdHPGSDlAZqFNy1UsgeoEI/hGutCF1XhDU6W7PWhblE1GtMIqqAUPcjXlTvOHN
0HkDizB2zDQeaWGC01Tr5l6iSXMXwTxUn/bPUv0zgveMAT2T3prj2WRARPoIu9KJ
dvlX5sw5Db8nRf/++T4GCEtnbl8HUNwh867nmdY24JbPeDemeoEg44I7X4rZZdcT
hnrmfL5VL8VGf2pHhT+fLYUkNciqEi9SpIRsqxZHZS+zpeg/3c3UeRMCmNa2IXS4
Wxf3acWHt/Nbe/7N/ZX5JHBQRnMrtMo7P4U6jhtTL5aSk1XAJXEMj38ehhuoeFRk
Bp2LFY5Qry8JyE0nVKmdOhRYv7+ddRpEZjmHLymBxmNMA8TWuf20/0dNCylw9zWh
xKtvLjRYg6rW3HHp4I0/ojdkxZueYat8JFuOffdaj2FaKyyHA9NaUTkrZIUem9pS
69RaskujDUZLabPnl6PURRZHxE8aUEW4gBDplhv5w2I8hV52tWp2TBtzyFhYQwLr
i9zPeEBhSanKSfgjGMmkQq9zoyYfUXVyPtE9kK+2+LgNJFl/cS2l3GtZJSbN6df2
CNILy5zoSW5276gtf7fQnwstI8IdwgKOYsLX2Dv6Dx6lbA26o5azUsLcW0y8LgqH
Sg55Gz3DrDezvMCQcTpPeNl2BgNO0mSO8M8t/cnpqDQEmcriBRtwiHwsKHDDihox
9rh3AELmScDtpW2eLhtK7TYmtuaZGM17iNZtgzDc+jU0Y0h+4ZrRFqh+7NDxJzkn
H6MZp4BiDZxDpY8Cdc0XNoud6EjwDj++WUIt2p960bFOeP400c1CBs522WSjE+LQ
dUo4TyVEhqgd6eaQMJS6GYyFTQSGjutuJUeSiEbrDSQYxUD2sOMZO2h80grLGidS
84edv4/s8rpC8Fy+YA3o5aWIby7lgNbQ9WyMwD+nSqtgrLJPyKiD6CqcK0IcJIY9
WUhgLnLQJlajK3JrSsc/LaHR1IuBCMERq1hkh4QSuC6SN83yDY/XUAroC5d94Qt7
cEZ+QusRlh0DKoJcCSGu13AGcELAZ/vFebTCSpIMKuDZj+zicYjZ1KDP4HIYLVeW
9ki8zk6ZWB5xGUZoR3wMLPKESyxma3AVFzUuJ00leOx3jcN7Z6XRNEYwiiDqhUfK
SyA621avw17kt4SeE1TTZwcINQw4b14Y88xMXwQY1qU8lAHnj3oQ8Ap3geMIglPz
SyM6pe8fmoZ9Z1mvPHJasd3lKKwzRRWW8LnDYEWDKS+JvSjv/xtob/rwNL1opR+1
iVvGmp24io+HGp5MkcYiNKjgibfZ3Trjyl2w+FIJcGYGWTb6lv3wck2R8Ng+lope
ae/SQ2TgKBrvXn0wlbmNdfDff3iJJy/8ymf6FxeRHrqMAHdMCaldkP6cQUHQl8Ju
r4dX/tWlUwpOVCFiJe8s05gqtAZ+aQYeNStX+YYqo7ryYeVxhlXsk+HB2TbsR5Ig
Ia4R8mllUE4ruIV18dERYAmqo7fjAcdELerJ0y9ygDdQveb3BOXkN3TNIEFiKM7P
T4if2YxVKY7vypmtohBAK9ONPzIcc6i7bjWoFX0itDK8T3cDkOBouLyYBb7fhhcK
dfCuaJ01LtGD+OsrvCaDeozpJ+wTvLKjFYo6sn0TakHns6/+95mwh3/YdjUA+cxR
D17Ndgtfp1MuLcDiZlIxdAz9Ke52XYAJmhI8JLiABAyhEB0nqY7Sk71bUGeKm8Iu
2BSJTviYCCTz++vP4sw3ZVJRQPUDAhtqXNd7rGB07blFPYnTPTy8cVHg66rsGrUV
E/erm2uCCo5N+3B6ROaTSkwGN2v2QTTyVUFKStkpRSNv0l6GI6BxHXdPDKHbdEqw
tdJZsUkYS/EuviCln0f3DAzaI47DO9UaBKWWCAgQFSjLKtt9RSrKE9isCYax1kqz
KKljPcFvgN3zgskAL8RFfSprfmx8IpZAMuNe5aUcJJVMNdnukAZR/0QTt4PYUuVU
G8adm6agjTQGSF4bAF4s8pqcM39Dxl/OYhH/eNbjAhIU5vQ9loGiFnn1bLPyNjkB
qRrwGmej2pnwG/5Qj2j8XCAEFzrn36EBu/rwpGANnc7YUyFP4hgsYTIuOnt0WAjU
88WxRHIJ+hhxk32lokh+G3U/+o3Rh7jQmiTzK7545jDyL412YYcFX1agL3U8aetW
vUVruX27Z6iE/4Xh7Vi5gEEHhkkKPQ7OD/d0eglI/jMpIveGkHQJHJprt/pQxUkM
DwhAv4REpNuUUoFEL6fKjky8c9j6emlnI8NhR4zlMPQxy+CCh4SvM3pbTokjb/Lb
MFUsW4aNfOLkkSb97fyLe+RGKY9p1cQV8VNJM88KgroHqaDbVMLf4B4Okm0Y/mR5
N91D66oAkfLELav8QVZWvuey/70Ejpnlu459xT5f9NBF/bGxvZD7siw4wbD3nMFJ
/++26TTnFl1ePd89egfDZPLV2st+SJn1SLc1xIhAfHWqjCKC2U1Fgy9m70C3xpmi
mCEjvAwG0Ved8FWPz5D2uBIW4XAka6hM4f56/JhSAdc8ZLAZmLoHefHsFLnY4UAG
KROHghcDYpP5jbSy6lKQGcNjzworQUyNPdBEwfEMncJUwvn7wImRZJ/mFdZ070d/
P0eQ1bgq3WvFbV7cnobjzpSl474jvx7nZh+wjePFZ8Kez+Py6Ma/fSTuawashPdK
fi2PZOAr9MqDbUP7hqix7dZbIQ6AMOu9P9d/uThdss3+/2ZEzQkyHBbnX4hAyal/
tVplFdQKapRvQeyR+mmSulxRt2zn+Ra/pp5ZzN0E+bj7zbgV3p7jcutQSsRrRmUj
qcQwlv55ClmUJc+MvJbmNkbTcLNChIsvx5KgH08LXey5PNMfpR+tiF99mFtYkLC2
JWutFqvpnhsz3kIWklUET0q0bRN+Vw5TyW4FdL83MHanb/btxRtFetb3v+Jjeuly
TFfqNcROyFHQJKwhOLJowQbyLRIMMnW5K24+g7N4ERbaonTJNLuKxu/hNQaX1jZx
CBjo5kFrhYsa1TwgKerN1Bi2/G98jSPKh3Jm6weR34sS7pBR/RaGLm3aF3nB0pxV
REq5UQ9gV+UyRo5Rezrh4g7SEh/USHuk3VSMVi6zIrvxgUDWY24a93i1moU4hwBI
mO52sFp2wKkcJcD4+ZK07GAYTO29+91JZIaMNTs0HF0U+rv0aunjgm9xprgW5P54
W+rbM728t9anzEgoUwmtPB68UcQNCD9Ps7wjXGoncpmXsxuhye+cPMcYICZxWwEE
2Xwap35rNwWmP920cNA/8LfLkak9s1Qs/rKwLqskvTeocT8lJ+c94I0SPrfwGXD0
ol32LKKGuzTprj7ZNMICSjOtbW71Q2dqhVa1W249BT9JIbnMigXgSbZ7OM5KH1O/
rHP1R04BzKhoiJ636fTz+7c4pdAGz4qoJfot4cUO0NlKjThsA0xcXVa9XbNcHJMc
iUCs9j18hA2O0ydiRzl0S79SuB42LA6EDmGKvC5Z3Zbxgr17QCQ0SHzhyE8J3ovo
br4e6KQpniU6qOmTFgEHrJ6aeaQdgPE0VwngeheG+hT7UJpWBl8sKhiMoZTYsfxU
bFXXn0BYjG3Kav6MTmEnyNkeWobhQWdj03jJLXenKVZWp1NqC9efAaUwwtLPi4De
7aMOd1kgmetXCmm4VrgY8kwtaWfIZJ5ftXNL1+92XMxIz18iFhqsglGyHMvmVDDK
43HerlZltgwTKm0i1fDPZ9HhhTI49z5erS8HdduzzSKVv8lX8EKdnGqoB2clcHDI
syeL5PbmEASyDvYWNfkdc0lbsguaYkkAWhI8EbGDmyBfMDZhluGDJ3rONsl9kNuI
`pragma protect end_protected

endmodule
