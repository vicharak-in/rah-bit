/* encode the mipi frame to send to processor */
module rah_encoder (
    input                                   clk,

    input [TOTAL_APPS-1:0]                  send_data,
    input [TOTAL_APPS-1:0]                  wr_clk,
    input [(TOTAL_APPS*DATA_WIDTH)-1:0]     wr_data,

    output [TOTAL_APPS-1:0]                 wr_fifo_full,
    output [TOTAL_APPS-1:0]                 wr_almost_fifo_full,
    output [TOTAL_APPS-1:0]                 wr_prog_fifo_full,

    output reg                              mipi_rst = 1,
    output                                  mipi_valid,
    output [DATA_WIDTH-1:0]                 mipi_data,
    output                                  hsync_patgen,
    output                                  vsync_patgen
);

`pragma protect begin_protected
`pragma protect version=1
`pragma protect encrypt_agent="ipecrypt"
`pragma protect encrypt_agent_info="IP Encrypter LLC, http://ipencrypter.com, Version: 23.7.0"
`pragma protect author="Vicharak"
`pragma protect author_info="Vicharak Computers Pvt Ltd"

`pragma protect key_keyowner="Efinix Inc."
`pragma protect key_keyname="EFX_K01"
`pragma protect key_method="rsa"
`pragma protect encoding=(enctype="base64", line_length=64, bytes=256)
`pragma protect key_block
KwFiPGsAmRHO5/MnYh54sdFVrJDqWcRkD6W9QDJ/bLOuWjhiYDTG5wL+s/cdQpBs
lAlN6WEZ/FuLdOgZsygbFkjYqT5gaGcN8LOMJXABwb2QBUeCB17qEc4bczSfqcjv
o9A8g/rXV3EAY2m1ThT5gHbzFsRW7ftKArctMQxm9R9K03ZmFQ0ayWeImL3HQDWB
SLx2NoAoRN07pbMRc7Mc4apEq2RlICDBG3acurKWlW4ZnkZoSoFdc/MhwvWHz84d
6tRtriUM985G2EfFksDkfEc0RraFK/8lj41ibBxVfU9s4T7em2qD/Y7VqZRG7C2Y
H60+AtjpqikMOzkEyQ79sw==

`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-1"
`pragma protect key_method="rsa"
`pragma protect encoding=(enctype="base64", line_length=64, bytes=128)
`pragma protect key_block
ZaGdDGY8bb2JQTlfNOMCnzjet4NWFk2Jk46gR0P658/BGeIlsZrwCF0FQoFE4OmW
q1RlhYZxcZVU2T/t/pKlF0epTp03JWWTQdgt9XYmSpWpGVl8m4mV8lXh93EROU8H
Lm/pRVqhYr9kDpr0e/bhBC344HoMZsHQizFzm6E1TlA=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype="base64", line_length=64, bytes=9662)
`pragma protect data_block
im2OdrvyO8cZcuzdT3gtSTJgjZRn33X2S5sRj5mXc9GWemiMJFtBdE57g5jvmEaa
IsUnjgYWaMEPloUDTAuDl+cPB/mC/5YKhpk9mCFc647qkG2aGWUNme5K5WjSx+OM
8Wb0CmE3/dGFI5+2Isz10WmhqDw1JwJCUj2uDA0wfqgdxRqRyxHF+ahzHlTTb0hR
kI7AssbeaiTAJogKc/GUdYEfXuRvwW43Mb7W0rfTnBsyQXse9YdsaouqlK/tnYsE
bnkWyqvmbF+UZlf11ZNJ9yvRTuDEYoUUlCDEAXdAtb4Tl1I1hcgO4pz7aeylGjmt
RlScRsT5SunTxJ6gBvTzLxtfkRDh24gqcOZT5FDxOrhUf8sShzj5fy6VmcpxcnDk
WECsyaBkFNycNtvjnAwKfE1BgSfSeTc3E8I7lEXAECOY5w1bz5B/subWrXmehRMx
2Q3uFiZJeOLik/wynnfbAHO5cYtNuOKQeKb9kIWcrfjeN3wFHW6KkDFPpyXaVhrz
Q/Mi/PcUCrNrQ3kGCRyOYCtcBTgvyIfyut9emDp2rfDtSVYAFb0bqDjdv0WToZF8
OMZPjEER1R0LY3lwqDEeUBLmobP6yVEbNQvXeZmIyKeRxwz94cMm58kkSwpC/34h
L4njanH+EE0CQLjwsBZ9mgnjEoR2/looqFFgaITqoc4y5mV3HkGuR2YigQozXSE/
AlGXLKorO3LRQkyG1RxrXVOX2QP7YauyUwmhnFqKNNR9ynOeDTazrsb2RHZLjKAz
90plo2YZWZbxEExDoYqvIpPJTr371XerE4e90RE/pqiNPA0610M09h/2fKeUBPR9
C0AN3jA+W+b5xBX7mlSoWIOAcLrGbY/sy6F6NgKYXAe+5Dh0Q9yUOJPThMZg2hXV
VPeNnrFY1wOuyD5VXUdde0ER1tng0BQKibMh9ms0BfyYJmyN/9LGO+cp+qTlqfgJ
2pkIXUggwdEr4kR7/8Fr4r394KRWP2A4GxmJtVK/axftbS59PWq6Qa/PUsqUJc9J
3zCHXv/FwTxVN4IM36/zG3ce24Gr5u9vifvGWceAGx/bZl3Lu1qQBNhNreJB/4W+
Uf4SrPTlFBUdgAlVJc6rV8Ef9H/V/DMozClIJ30zf9cd3hazZ/hITTZbdBjEznui
n+rg3tJHG7QuaMjYqhZKDx3wSnyD0DHE77Wk1pFmTBekl0QabbFpqA3JrRVlTGLD
xVvaxuT1CtxHyHAf8dzLuMvBHjCz81ewMy1se4/JROhDWwPqAMeSTkqQTIF1AXQE
UOIi8pFa79EcaVpDNQ91TxP6IeZVM5EkFrepjVTTBnkvMtgd0e2lXzLbxLMAkDMx
chOdiA93f/futPWKhVmroget2CwzHOfb+kjfz+wDIgkzhB23FoMU0Ie4f0GvKwXI
M123e4D58P/GtrZo/BU0GiEdUXiymY809Jvkp3O0LjJZ3FHAYJ9HGuPVVMD1dPGf
o++RrBqwwcj8tcVF/TaefAYm1bcAr+HyZKrxCGalHAPTMNvCBzeDZsvVAywwKEF1
w4Wt9x69N4YY3XsDLwGv9UmfBe9UaZ5SkWEt7ebec+PggkW/y598dlQm2/2Ikm4A
JONxNSTrEdQaSn4ewQ86qUGFwGAJ4VdxkfZuda2UEgFGul7dgl+wufhZR4R5yr09
WrCB9ICmVrIZUdZ3fLhOk1R+yc3yMXwMZLWGF6qx8ESz2qnjY+A+16CJulCl5Guk
N3xxHT1kYHu4ItPXq/EpcvkpPAAG1XjLoRW+IAsXFMeYzDYs6vPVuNeJo7yTZAyM
zTkVWVSR/K3SuCJEkzfzQqWES6BFSFBfY1aY1KnUHEq97HsGLGv5fbxNSASw+DPE
s2CZ1xDpu4raMK0TCl82SUzBvdjFzK5U5dZOXElMxTge9U56Q6r8FLK/l7iTIEyq
JB1YhHZJ3DHNWmmrOaWJdXZPNkEzEiR1c7wgw/bl4rMPhgGe/fW0m19ovTHDVJKr
NWGtftajCg83UEZkBqYGNO8SR1ypFoMX+EFs8YxU504uCcLucgeUMswkpOW3PS1A
E7IVKYx06iWAbtdRrm2bcyW/MYUwXTasN1YS31w46tmuFA3B8OyYrc48ysrmt7uM
l4TB2Qh9MHDRXuoOFE+m1z8fiAnotrTQsP/4pnyGoaq7IGSx3Sf1uOF/bem1Q1oz
etR0+K9Z4yRm3OmkTftq/vRakB4r3Y8c5MOj+MBBlFH+THcuOgZwpN/vuei1ZezM
2oZ/iU+XxGec6JH5gA4hay9Wwv9LfzTTNxvOGxSl7os+wPMAc36SfTFsZ0zu5T4m
vvjHt0oi6U3ESSz8JsaP8VdkQqANCSK2EdHLC+YGh1eizYIj90rD1sbjoQvRrGve
hKRQCH0glrsWxcmSMFO80VTQClOU9adDGc/lsSIGoI66QM6oYB8VKESY1XWvW0FB
kg+O2WOeGvFXhgJic6sOwSWJmJ6nrNT4zgvof2ecYOU65NANAZA5DXqsKXxDIIzK
uS7QJPjRV7ghFjTdeTpDGDZYzkNKeR3yDrXlwmUnektxnzlIB+olAOquH+pPCN3b
HFd5Q2q5gmiMzFBBTTPcmb7gKHnxzkUxP0NGsn5Ho4zg8eqbb1VC6KhWMYCsJ/uJ
4xURa05kXusxGOk6innWj/fQFyv6KoMg83J69RPJ0IV64ThRRls3giDvhcTtjELx
PCvNwwktpWwpG+m605saWEIVeQ95ATzerjxmeM0q/wBNFaeiIhp5uWoAljBVh3NR
rGIz7Lq/LY6OJT/fh4MKRqxd/MhsLtDxfFsrgLrezOgLLWV0HetusS+Pu4Uoj260
bnwL6CHGKIZ6YsPlt3aXwQtcCTypGtilO2qpHnqFG05SinhQUjuS+fN8mwWwJkyx
ndS3lHPOC/ohDlHrGjJAyN4gSeL0kK/nGqt+Ni+HP7rWeL1TIpPG2sP8/5x4hpqe
AqzE/zIgxodVqV8Ei3qQufquVJKWMTtRMS81VkxVuwfmfcEE+XIkBjWiiak4TxaN
ZbbvOCTqIR+2mqxEdyJeQmwVflYZkLDyBZuPoVoN8W29MrASCOQHVQT1pIw3h99x
HFTdWGddgShoH1VX/HoFzYK5SGY/5yrYeSuPLl2EGqShNU29rrNYTpvX+seFlrCG
hK0NHj3XvmtvHeDWjDZrNJBhuUI9TpPfZMHKy6VBcXOnxj9z0qhUo9Ly7kI1uT06
7hJFtwVwi2ncVGJpZy8c30tBd0scF+KOuljx5rYmR9PAySdaII8UJ1oARbWcufkR
17oMp/eRk0w7SnTSF986CokGjoCs6J/UPDpUKzdn7pCmzfIC5IwkAWAFpgBzwL/s
pr4l7f56e22PU2+DeMX4XekdVvZTImjcm/pwvLCZ0AlGTCz/t2RNh5RHxIvj5vrN
aeycD1N7acp2M1lBmJHtaZ99fFOsYpoFgGPm6L1NSRzhZUl61GT0cmYv+mm5BVif
J+ePJOAdYSushavOw4PHQqIc08zPQVWwZE2hHrH1EwlkuaD+37WF1TeTkZvQbh5g
mQIqaZEfzLeq5vb5ymhTs8RhxnrLfaS2sEEgqSQACqPo2KnqnpDLSCrROe9qCYFP
AJjwdDZlQnwxDBpXskvbutEuDbuKO/M1wsJVu1/ppRgb2WoPfjhDZ2pZDxGaUa0z
m0VAxp34G5oPTAKScaew3y8HkKivVek5r454r4BKWxP3jytTzENsfOh5L3vbQ9J9
dqOubMs2Wp0gYd4cRjdbY7FlWoJooXDKKIEeV3m7c3ESHme7Phg1MHZlPx041YhG
5Im5q7N7cH2V8APcE8TqXGHIuBts4vlBnAhMRLr7FS7C5X0unIWOaMtmyxyPZQPk
rSTlZtPyA19e+6f49uQIjc2tzyfEUJFrOOa+8djkEVmYm3CEFFID1ULuogZLPdJS
Q4rintZ38t3EV2sf1WAyFkcBmiwQu3kAvtTspBZ/R8B4/GuqDvhRDTFEPru8wuMM
jJvEnwSkZ61ktTOSVYXqxIm7bBaQOXZ7vWpDgi/fT3d5CPhIDBtAjDP6Ac88YC9D
9JEaoI5zZaD6xvYBi7DJvfxatXEXYDp2iTpy28U+VDElBVjRHsIGwKcIIUeeTlqj
/0ZhruIt5yK8Km1OKxD11wniGpNv4RUeXIibHVhDq7K7+OfA7CDrQVI7IukCnb63
3U76bHt+7XQtBHX92+Ez8NCCb3qpJ1QAiH1QGVDWT6Xv6GJU/0Ik2FUm40yaKwVt
6rZcZTII4RRV7G4PLItJEJclym/ej3RM0QVYvjyHBRaszm7eyK6q2T2l1DpxaYnt
yKcxJdRDZP7CFOZPcosAoySj0VOiV+sfpsqdK+SobqYyYJzda92/M/P+D4q9GUMF
m63mkQBomlm6nbe6OSmykDExuNTBEf5yq+KZOouUZyD9tYgKVJ+w94c1HXP7cIsO
PZ68V+hWMyRvZM2gQVuMGPLMuDP3c3Yd1sttaKkW3VOlkFl7wLIiQg9HM6Zby+iX
eKW7op8pUhFUkdI6k4o7rti+b/o+u9wmO5cGexkDvvvXbkYwGEYEZgyOuj6BUiCJ
6i0FSuvG8tcQ+NpxWJmyBppbJehp7GEFGr8MZGQAsHWEbUc3WHnMsM0DAUwR+9Qn
TO4lXb0YDk9Y6XTQAxFxYXbehSJjjZ1QWjWalO/5Frs67+KGjFCPN1azhs3mCZ8Z
otvstm/9RyuEzV5rEz0j+LOlArsg2TRvpTJt6XnW4y724OdTai0UQOoOXXyPvQov
WU5XdbVCse3i9Zy0d3OkMDvhPThW2ScOETvoO5tpIfjjSgUs9Hgy/8POpJzGU/rG
3P7RNyFh8cEBZH+BIFcYOPor4mJTnEX6nQSEA1i0y7978wtj4dcEB0be2cVaBKJY
YW3dCeuhBoqD3JDtXCr8pPrdbKCuEwf2jRoC1uCiktMGp7TMT//infSWiWdnCAoS
7KMqDKoDDsZCv3h/7HRzrwRMV4LVfxqL5oiDy4wZfQpx/ftQ6NIZbvt1yXPY9p4U
PUaUq48W+xamUnAXjNCwkWDWntYpib4bVZfuRv343YIWApD3CZ9Q/vePsxsNfhfg
6b2LF/aCkgQlSsI2C2oPAZoA9uCx4ZPgVTPHqeXi5ImYy1VUNzS82zs4McosSflE
NiN7ztwDWYoDj8+A0AkRlZ/jmEAbpwaddnehIH2PYRq+Q3dne23NhHdcpIvbnX6X
oRHhMAreER9Bh5FiRMKSwzbMQlZ2avdsUK5KP5l4UX6fOX1mTIQDicOIXSlN6aUs
F5/phXaMlsL4uzG5wfcqNpU6afAEebWQ9T5/6wl+lTz0LTuGlUKJXBCPZXJgzhZ9
epVMTNVkxvBZb+hAMzAJQJsN/H7WMkgx0lOGocFHzvvsxMCE5K+8M6Rkv0m5sw0+
mnLU5+zISP1KOpSjBhJLwgzoxbBRo4PM5rU9a7IlVUMh7fjADA6gg6lm1x4DAw82
V/AL48576GVlt7xRjvaPMLBIKWRm3mYqR5CLNUEpO6DnOTN63rxkDHtG/JEsIPLX
86yB+Ttx73TkH2Fd8A1WcjMjXiqFzpGVXfoLgJb3ll133xFYz9sAnRLpJQ6gdn5E
yYa5PYSxQNNVJbRySwHZ1Oxy7p4TetKTGXyQryFk2NFN6dSdJcCwED30sKH/xS+C
oi020+Lw5Q1c1Re2IDwnUOF4XWL83Gii7QBGHlXN4umXydMda9X8LMdLSHIIBOfm
ggm2pfL+lHkq2CYYiCnm3r85/1VOiViEW8IAg+GYjnS2q0AQsSgNGjzERPNijlIX
DWH3n+ocM9MxHYlOkRXWOUxhio+eSjVy/KyZ06GlzXCmIwNg9M6z8AdcHU6Xnzrr
e8EPdSnFhgEwt/ZzBjWTgU3PGw7C1gDjU/068W6KedNafmQ+hZt9iTzyiHnXVXrn
UPgydla2V+eq9S1/c6FLiJRtPYGNUtvmYqzjDVCA4wyqsCNdbyytqbtFYgzaAmPT
uXCfmpPrlKBFb9cW/DtQAtg4zLgWMoqSDhs7qITyZAyu7rIviU6wYnOPnYEIWj7v
4JlNMTIOdo23tSwxj0zwJkbeO0eVgcixar7DadqYIrbPyISw4X5nBpJXoOXQrCxt
3d91a/RPs47E6OdSU7np4Fv8C/HuX/JmS4yTRxwilsntpTXk9obMAI3+2mIwVlJV
8tE7/CF8bStMFCQq4YmSU9k3UJYk0TsD2FveRhiOBJe1SwoP6GiM2B+h8oekyyCx
C344WkcvrDtTVM2r/qwEMUfWm9yDLaCNHoj6JZKKSqkJ291MqyCbEB/QIu2qO/lC
3j5V9CrOWDUCBp7WTGxZ/x0mSnbglG/brQN1iVXVhrS9X9d1l75mZgKiNIplnuI8
5SaCz8hwcfRCoUVy5/fawoYJS2p++xn/pMTV2pL6O1PJgwdbg5Ytpd5fpTbQMXhg
CK5omExYOB/CmFVUC4PALfdn2eC2csly8ijBK1JYg4PwhZ4hL9zZ/ddFfOKAulxC
jntZ9Jz0CJORj/7Xn1Swdasno+L041SFgmZ9Y6qfVP3qUfzBM8ETht+Mo/knt6Ah
gaRz9fbCwS7Gux7ZQSfKrRiLJrd3l+tRBgIK3HcXRBwrGtf5MM/T8qZt24Ybd3UH
F3UdHK8bC0Mxe7vzzGHew8dp8tdgOYQHmmcUTA+R+mNg11N63+ToF3jQzXG5/fO5
qPedEUNhLiCWAm6FPhLCiG5STGaYv7Wc1RJAGG6D892lTQnu0FZciyty5/4ukGih
MpHTJLHzP3FdPOhM9rzC7dTEqMIL77WIBuX4gtoLp3wf6VN2bzgGuWL1+/WNSVMK
PsC2fkKgb1l0CrdP+qKhPVxxeM0ADeyaUluATTVLhpzdrGJqDy+2oPn9afu3pOdL
PGEA9Wo9+HBvCCc6QKN7wbma3h9fonZWhZp/0BPtB4ePQDnnTDKjYF+DLKVit9D2
/Q8r20F7jwER9uH/5V/IS56wrzwMVGY9Zo4zR1zboigPS1fbIf8A0UUdfekTh+hF
Z+h/K6wseMQD41bOPcZm+FldSBGzhRTnkcCRnW04ebaxy0AJVVSnw1rvVevo7Esd
Ay5ke1u0VgkPdWNerZaZNVUAuezon8NcNBs4klbrgktSlAij64T7YzLuE25xfMk/
pb2i7igLRUeUoyLNgcqYXzuL5UsNk7xx/R2+KOd/5vSrBEmvr/8QXGMuzZn8/RwD
YXVL++mbV/EZkvV8mfrqdMFQYZdWf/0DxXtkwiLoaJL7HwG0jKdZr7WTDKe28cgh
8YZskd9vvjI32hX6rMFpiE8nWST+vjYVQhsdsvkjEHwXYOPnxZKMywJTv130cSDt
YpDPn/nH18rRDiEv50OHZb923tGuXU7KJQEry8BTnompcWIsBwTv8+FOCME2xE5I
dUMWYez/AVo+2Kd4avb2NwPVqWhrgXgnX/B/ka1usx/dWGlIw2qBVK35OgKjgmgF
+qs8vhyYW6et72MqZjqq+BR5T47mtv0lZzfsRIVJ5n8zDRFcMs+ADObVPL0HUq0f
lwUOn1RzGTKKGbtAcDoPGJlN4rhaSpqn3LexgR7hifyWPUmC/64OpA8NNT/QxKC4
rms0WOZotqY6Wq8ZOVyfVlDeiOlP4kOXRVSPOGfjK8tHz/LlD+L1kFj0YwXR/Fcb
zzOEPGY7UgER5ualzatc/R5uy36J6osy56kyEYp7PL6PTHfSpbqzQVouuGKHhg7H
uZHKE6w+9qKIIhgD9nWRl652/rnJYIorRpzHImVvhNdbX2C8bKHmE5EKq9sJvOgn
zn5xFYubyCMsCA0/5rLGynZqgfLT7igEvTVm17s+Gaii+6szGOI2imTa7qu85Kvy
DiSQUvXOYYBjKXQAV0uMoajbiQrFy7vH/oqElvHkGzUiwNoxX8O2E7xKTzzrNAeu
H1k8zt05VhbgTMOwFka4JJOPNx/g3/dRMrrVeiU5EE/NDGPJ5gbNRbjnWLiHNQTi
VojQ7ueqXA8diq76/RdAlCgxJJ5hi51iyorvMuwkda3yVUmSDp4cQn+wlXwo3tyP
iJAyrFuQJCBPA8OcNv0B/7KQYbr94YDhQ8X1XjNpTHtuebPlkgQrS91gMaR110I2
q1ggOtJOG4qsa6MVg8BDzChr2yv5QDM8EZdHiM2lB8cQI3/WMNgiUvx0jAn+paDd
4ewwiEjsxVPGGWvSC1dNaGVp80BjaFLcgsKvW5JY/R3GGa/d4mBUzrsfTzO7oS6f
Al68pTAvJGKLC7bG8QRNTAQSDJp77sj9ufSKBEzKFfbK4sKJSfaO72fqt+2XA4hQ
one/jzadPtBloJisGFTOw7qKVDe5q2wBtEcbL0hCDwfV6lS060/ApKLkqhvRfqrN
vJgsAGWgpa2wXcY/nzfLWfufcPYUyXqz+Oo5vLCMCePzywsx8Xz/Q/4FHHWkZfaE
NNwMQAKjoVJQFIs+vIiUYnYsEHioUXUcsDVpoXg1VeNZv4Y2fyMJqPeOdmawk3Jd
/TFZ7p/3XoOV6wDfLEoOF3M0Ttzm5lCTeS+5EXYYdjLtp1Riwbv1PbxDUth2Vq6K
pJHumW+l8FpnbC+wYDyuwrHe0Grz8gan5LAPmpZCfdIV9l1MRzvhakVc5S+5Ky5g
h7AfMYmZtlG4xmdVXRAzKzCNsHzvLbzcoLksy0/rNOMtOIo04F5hvY8huHCTYUOI
ofs5rvTjcBLzmsi6BgVerehQ0pLeEYGgPgL7/RpOalCrOiVYvaw5GBoYsQcDCUln
P6tV97JSFy9hag7Fnl86ErieW01xjrKA61LjVVH7LcTJl9PJ9imkN4EW0lzXbXvo
59n8aHnzhOMTDs0GKvNpwangy07eO6Ki+/Q9Cv56fT45TmDjlS234TeO0AHQnyhH
1dXF6wHRTC+YaiS4hGjCBg/JWhgtUqhnX7hoQpojpECFpkp2D/kJUxpX+ldGUDsS
koWdKWBe/IbQDaNGtDYaVs0wz9WYGBNeXAfOX5RD18RYvFRs5rm6PjmQvKZPgw2O
HMsEoxSKaJ+P2QVhHTfL4mdXuJVgrqjh5WfcyU8kiytO4gcjz0u+9BDJtOVthPkl
MTML3CDBCtM+v4NEyqTSaZxYSloUA19ofA70XbwG6d3L+qPUq+tydfqTWnILpHky
egqg4heJ0jhoWwcWbCdxwjUdZ9xp6q1PN5yCJlW/PvfdeadjRm0uTFctTJvZBzH0
9qEtq8N2y8ALgmoP9MxS9Wmc3mz7j1An7ye+EL4TgeOLpkfyeB7Ug8Qy4Z2pDFE/
C+yewzBuZKqbdSbpCPt4uLFRrphuxYmes3rQTlktDYYWyvX7YyL8jiJnltpK/Lr0
8J3UtHF62S/l6/mRzD0bCw5qJH5XsyY+khzakRlVffE0VcSjv4t0Y1hgR6wZtuT8
8HOXxveZ9zf33apat/XXBQ02E2HbY9mHQLMZHNBwC1lhamir0kJtawDCABrd9aAZ
AitCEscBp8oYUFxFhXRdwCeqx+myh4NfwRuu2S9F2YPIyIvOCDHLFfl8LCoP2gZY
Urpg9H8SH3qKYs/E559RYuaQUX42UBsQehQ9ST/kJ18xw2UQnW2230KRgKMqzvGG
4DJgBAhwnSZEuASAG97sihY5icv98O/rokfuh3tBwedCUlXwL1MRCb9+H8TUJDM2
iaJ4BH0VVJA65bSy86/1oZK34QIF2zIyBlT9f4s7pjahJzatovrD0wqVMBXFBvXs
fhCmdvhTyQGdiCNXva2xwSAo69/VP0mvhSwmG9AqveR1pv8U47FjAvBiVr2rfKSw
U+iMkL5y8iDCJ+w6/YsBIsmRctW3zLpobjEilfGtw+BBebuRrNPSv9niH7CSt8v1
GE/fTs5wxvohfoExC+zVvK/+dgYYE9byOc/lv/qpJJFFOxGpAWcgF1bx1KBxkquY
MuDxTlPI0XBLw+W3HVyGO0Ts6B9vfBHJQ19Brj00E0dvK1BO59+2FEA3TKP9fN+B
YeKsm8OTteKktqOMInX2BlAIFoOtmULGJddoH7Hisc4H3PnvweLcZ6mKOCUldVPa
WBCHQrFNmWbUlMBeDi3sNeYe0ayoNAVLt5cdqKsZahYdJg6R8w/gLJU+DL1Kwuj+
4mwTjtrlF4jkLNizMlm/U/SOkKqwohe8+XCtbspcDggq4f0q4YGuI2wMxXwDmfE5
W2UTPtl6ERqjO0fEpBZpnGqUxeXzUXXCtTutWt/IVYsWdUff3dyHnzb+cNrbQvdi
j/vc/edskA1lndGfS5PaXPXknHFdz84ONgRVTJUbpiCZaqLOPKX3vZTcMlDILDUZ
M2BvNlA/6RwSlNx54gjTbSb8OBac0SChcl9CU1BOj6lfYdQexGYq2ZZ129MUXEMf
S7+Tg1qZspqbrM99yYBfnkF9MJUoVOyOzSNzKKb6f9VyJ1RM04r8bH8nGXr6aF7+
QkDGXhJQXaX9eKBwPXLXE/+NQReTCNH5DWjNV5Tf0cCnkJeOp8DX1Fs3ZS4PEpHG
EHEGpJ3K4jeI/1YoLAUcCRAd7U0RqgAkUVVAZUkd7dAvzvKeqSrJKWZjc/TF6ntN
Fyak8yggCLmMgJAsrXVGjUamJpkjYKZRrEVh5KrsUhgdtkGe8QbdON+vZpECpxL5
fN2hg8idtKMUSL8X4bFx3FEXaTqZNXMDoohWjC5J0V+3ZfT+gB/oIm0uZ+lEpNd/
IuoG8kVW7eydnkXHQIhwy/phkQzKCA1V4cD2SKImLR7ZxXMmEwqxZfcF7usRl32b
+1nHZA/2MBaojiU33X4ZFfFXrgD/dVkqNZt6yrL6peXyt8ebt0lidw1wAuE/SVVN
u9fOcjWRFFokHXM5gi+Lp0ip+usOHizfDuxQAzHby5IxZ6RpP0daFfT60PKbt3a/
1+K2tuE+Cr1c6CE/rwiuCev6XzQF8yzm68OixcA7ku+ts19Tj4x+T8j/hRrbDiGy
m6uKJwoWaz9Tjp8oeIFR8//XLw15TYNE4i9S8Eh4RUuoO335LtDWDBizuAUew5Pd
KMbY/BVgKZs+pR4tdCCY9wy9Pb/MCSUpWOMqek61iSWKJLhpgKVCmZmg114NTTWp
UySzy2LIObYKLl/tdAhFyGcN8yzBIS1WHToxLoGwHp0Pi7v+lbb2HzWRgoGt37C9
EsMiCqxj8cS3vcE6+cPMTH333vHAtjmiNB5Zob8Oo38BVg9ZhSom2kk1mPhIa508
K77BCjGP/EMWwW5dE0zxzruaJa6cM8AtfhrdMvdsOcRTuTqVp5M1AhXCYxIF0kJ4
96ridrWyTcp0u+jBKpl2cqYOu5qPfoVzTDmynhn7ADokSvp2wU796voKQtIFedMo
/yRIUCtJA8fd/ukPdg1BQa2KJ6s7r8Ei1fhPSVHwHwgaCS3czWmGYltAvgv6R1MX
EqeY6RToj9ba0d4JCW830GcwG/+k/Zi8NXP1GSPL9529HSoDop97yIg8WjQvgOER
WAXjn6GFKcw5500Cq9+x1wBMZ40U2QkazEvxHN2Zx2xxPuRSdHq8pfHZnDE3DjIG
chJzkoHOsNCWAT/2NSru492K3uMO+RFy4mqEMKblYooLeYdkK/FsB82ns1JZ/O8f
Q1j5pB+3RdLdmTksoPMwZyCcufpF7EeP1riRsv0JQXTl8LtB+Pw4ykKonale+5Yh
vNHgszl22dkNYerj6A7/TZHhiSvQrnQZa4STinxyyI1SWjKWSwK6nE369bWhpliD
/DaLZwa9jhnXMKCw7hjH0XRBlV11tmWe7yhyLTW3Z7ExaaU9/L6gPFysNp5Z5KlF
dSkF64t+YSlD/EMs4LW7ObvKqkpBoFUA1EvYsOmArcaLjbMGaf5UhlJQ1179KOwA
bRoQoQUHSc08DZSyr6kJ+9hElzr9exMtBglLjScnz/Ls0qhruSQ3MsIQYnLPafFP
gefRl0JZsJuK6PmBpF/ml4zoIWxZB5sIPejTHHGIyB81lM3k/uI4LO57sKYYyrk1
IFjkFe4IHLKejJOgkyJoVUazcj+kJwybTJ6nhZicCjE6DUt1K2w3qfmnnpfQMMYg
B3RlBnC+sp1DhuDVKLkPw3WRMs1XqwOeWHrT8UpoJj1zwmOjzhMKvLWqrBy76scS
OuTSdk2yqtQWiAk7OadQsPzyTS5KsI4ji9pBSt1XHeVEgHBkIdCdJ+n3lK1UtgcL
0ZjLX5FP0Wr0M2WM/CTYD2mxNff1M0DQ/eqrno8iKsvDzrWErKf25j+GEnC5srkV
WrpRqenpT/9eBWx9QP3WfR2hv1FuMQL8npoApf3S02NrgIogS8sSNTASd4OAMsSP
83d6D3C34qOestAdpX4xg0qt8TwBgnCf3FfFBfBwgdJy7LZxX5hHkwoPNUZezn2a
zY/CFIT9FQWUDD2QqxWRZ7vd2X+W/5wBj/5/BnGuI8i0twM+pjRF31ed2fFjnYcW
tJd7+jKC36O3a49VBWffLmXrrfZmsXD7l1kenAjy7DzY1Tk9qXfaz0vc9q8uica4
MGosndEMUoywvvVYGtCvVFaZUP7zvK/ckrufbyT5kaSjqaXQ9yJAJKptSsTQZanh
1OkQ2aa4NfE2YxF91L37P3xMtfwVc58XvN/u+RO05VLED8mn6LnCabOM2Ixwe+ji
+V+JjSKgNfQcmvMZRe2/i34KqCa3i0Hi4isj7hM+9Z2Cvvsjw+jR93eotp2RLrx9
z9Fglh2AUk9Lu0LDZY19lWt3qFyLYZ3wSJpYDPnXq+NHdKcQgXJqUGAmJqvURpXS
aNjYj+btkoMUNUYTGTk4OHyi8g7vZp/1nDQQiFsKGrz1fC1vWlDshGVWlfulXJvb
V9z18FUpfTgMcrPtNaSRXbxR77YM7QCLEjpZ5PE9YW/b1w9ELjF0V3D31heNH24p
k/EvWdn8OLfvea2azfzxt5OLpReRoK0vvhk5Dueos5qeooMUMfK9LxIsMifCTsYa
p+kM5yAQLy3H3FdMBQHLow==
`pragma protect end_protected

endmodule
