/* encode the mipi frame to send to processor */
module rah_encoder (
    input                                   clk,
    input                                   vid_gen_clk,

    input [TOTAL_APPS-1:0]                  send_data,
    input [TOTAL_APPS-1:0]                  wr_clk,
    input [(TOTAL_APPS*DATA_WIDTH)-1:0]     wr_data,

    output [TOTAL_APPS-1:0]                 wr_fifo_full,
    output [TOTAL_APPS-1:0]                 wr_almost_fifo_full,
    output [TOTAL_APPS-1:0]                 wr_prog_fifo_full,

    output reg                              mipi_rst = 1,
    output                                  mipi_valid,
    output [DATA_WIDTH-1:0]                 mipi_data,
    output                                  hsync_patgen,
    output                                  vsync_patgen
);

`pragma protect begin_protected
`pragma protect version=1
`pragma protect encrypt_agent="ipecrypt"
`pragma protect encrypt_agent_info="IP Encrypter LLC, http://ipencrypter.com, Version: 23.7.0"
`pragma protect author="Vicharak"
`pragma protect author_info="Vicharak Computers Pvt Ltd"

`pragma protect key_keyowner="Efinix Inc."
`pragma protect key_keyname="EFX_K01"
`pragma protect key_method="rsa"
`pragma protect encoding=(enctype="base64", line_length=64, bytes=256)
`pragma protect key_block
kZVgat5cQ4/bqYEy9ht8kdRttR+DBInCFutiyWql/cPlJdb67P53Jc8eOHQPrMNy
6hTxWpCkR53wRnhLukiWJs6DOGmrKyn5B54tGSv6BjjlSd3uu513wksp4xULKnm7
mPlfUH/U+nXoeYUnMJ1vq0BhUy5Xrg6zemx8MlR69x2F8fbBzDBhqCNQ3ngymA3c
6TAcA351alH7LJNA7rsXpwxjuS6XOuf5NnZZkvW7rQkDNyjEMaWn7t1ohYypyZAY
JjIqWctCXwCd9G5V3+giYeL4vOmwFiwiyDtcsb47mfSxSBUnDy2dhx1CBHWXnZ4l
WvWV0mJZO5DxEoBxdRe+0g==

`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-1"
`pragma protect key_method="rsa"
`pragma protect encoding=(enctype="base64", line_length=64, bytes=128)
`pragma protect key_block
G0StUPF0yzLX3V5eYXrs4kq0oNGzGtNPAzTeOoWaFh5tsZn1RLMPRbzSq3MIlmtP
cjpdWgOpIJBU/bTj/tLPGOZ4tPIEvajhzgTqVZucyWIZ8nqnQ45aHpdQdhh6ydu9
A40bSUaME3/sw+ZFP3R2uj5IGQ/TCXVtiQo4tLYybsE=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype="base64", line_length=64, bytes=9636)
`pragma protect data_block
nAbR9vbXKcHsuu5lj94sNGhl3XHYVGUjZ3lVWjAhiMAvp2IeZOxN0UKuc8C0MS5V
zvp72ZhEux4JLo4TzFqrI4WSidg5TPszTLfHwFIdUQF24305hBEnCYglJo9d+Gu9
60IxkA5dXvTuM9D2xhLWXTriathTLobl7enW/qnY5mZGt7MF2PQdFqnUffgp0Vk+
iF1HOSux3X+GBnEbZSO9oPURIvwvhV55ZloE/MXJbFbJv99N53p1i+tzm6az59tu
6zuZ0PXFImKgX8Bdz4A5byXYdJWY1HpQ7QQMcE313WpFFHk0e9Cg46MSpaIi7x9k
uG4cWG1vsSdrjeixoSlQj+i5ySajiTJUXfMiDyIDWfEWykjE99IF6ukOUfnkfVdc
YnfvO5cj8o2oTyu0chfOcJ7rXs8FbdO8oiXYDekkVqbRpemguGqD+YoVjeNO8kOJ
wynE8l8FOmFpEOTw+n6xIkq4j9V/qfs3M4CKWP6CaY4xZsTeCNzrbiM8O22Td5ca
OHtDYdt/J+rMIUDJYqZJcLwomFh0H4Chmpe0YKJuhEgdqgzl+A9sa6s6XUlt/dSc
bNpPx/fD5pnZkNFd7dKEO/x4aueFmxjR3l7prNYpTjujXSZE6pM0thwK5JSRLTgO
ut85SDzPGhS4fy3BI4MLIGOOYIBTlitt5YgLVf0okOUGAGCe7Ole44YuubwwItxN
byeqoQ7u7lTlN7f0BIfBBn1AKnnp7y0hv1lpwfj6bnEGgy9nx/KYgPCQQa/p0uAm
+eYxLHzM6AgKEn5uCv/in8niYaU5x9Ym0+0PO37cjneR3AqJHJM4jnqLbR6r1fVG
qddd7Pv6A0fZ5UZB9ETSYf2LOAYhBA9WTMtP/fXFrWMphKI9woR0kzMV7JjRze8s
w/lixGrywCr05SuBl0KcuKVmCHnfcnE09u47j4KGdejSiISKlu6y2Dg+G87xwBcU
5ldE/+dGmnBfRdyBb4g3+XHn95Nzz2gJ1CDLa9whoE7DznfNO2r/HhAt2EA/zn0T
7+kEUU8SyzhEnNb5ifTHxEIwMeQPwbI0wuPqqi3h3rl0MmvgKd2+RTKpiryh3IAm
d50kvd4K6ylLmwROdEZ/sS0rWGgEZCBXF+x4EpvP1pYbwMUaOe0HEPlKh6I8oN5Q
JTCcr4syV46PfTmfiEm/DSb4OqKn/82Nh9FcEkBzqSFYDRrMk7fYAwJiN4doN/cn
F3EWfoVc7uE7UxezYMoCVNPi0F4OoqyeBAgDqfrDKGm87XsswRDlGNsK2wDEd+i0
PLLcLCGlT29I9S7FORMT+sMtcNgfGLgiOyT/YBIpNpNULz+roD++S2fLXTwhLYHK
KRR3wYFhdBHTLfqGtZ3Gq3fIK5xW9ES7xxXgx9NfGAUjJQ5A9omRjdw0uksq7Knn
acMm1i2jHiJ9T2kcMrihcyyawkg7KF866HYs4Nsg2OsK3yZoQOgWjUCwO6eBK2uC
iWPF57B8K78faM1W7juEEJq1Iwauzo+pCamu6MMb5eVOADh7RQV5w8utTExK416u
o6inRbH0VORj8X3ZiYpmYenyi7oksUTzPZ1Os3G5RG6NL+8P14ohX+3RFefKfVVq
NHQf9lOOWvs3yxUhRBaszuwO9fatnTm/rog826PKjprTgbwnmeM+nafC2sPksPPm
+oDYSWmiNgJ8dTdh677f8monPH8e4zy2NTz+8rnpth/rc5yQy+vS2Jo3M6bC+Ztf
cHt9kmNIP/KI1M+reB75skmE9UVRs7Lv2zEO0oPxCmxpEhxT3Iq+oYV92oWT23cQ
QDPUNYeEC2UuYKeurffFSNilbbvtARS8cYZlyA3CJO5AJ2ek5joNZaa8qTluljWI
1lpYxMzvQI4qx4UZRN+vcMEdibBNNHJQAb+U7S8ioLKRdXlBXLbzqfKxBLUJ+V4U
EXXqJCmazoZRnujKjMV80Eb37kzZKPbffbdix4XdpYVNDkkEdQRIv91lAFQWI2pW
LFbl9UenbupA6qPPxZelCpdfU7OwQHxa4RvYQVKEs3ANOXdrSAc/c1yqJ4z6aAfd
xe65k2odp+mDmQLa+3LwQWtezdA0QW/T06dnpI7mWMvccpM3JkxJl+REGqZAPECk
gidekyRat5tpUFDxxGpBa3vXSokymBDacmJjPi0zfRmxY5mravNJnHya7wa8b0w7
i12soKN6OqgDRP1HxzAzVM0Vf9L16jzqWBev4xHjIJUL+LfGJM5L0hE5CR+bmOti
SnO7ilbmKe7SZPRxW4hRvXSPce9zzlZeM5HwzmV7Az0PCfGQBVAUGKZ0fH+EtHk6
z1sExYUnPPVGdVdQcA+scqpzMHLqnNp/5n0MFoiNCpD+Vmu8CaMjXUnwh29nLPLW
+aWpRtqg9KeDoDft5O3Cr9sxjbrwTuj25AsGMooP10mxle/TsHYx0zKhs93JHJST
34ncxxvGD0s76m5IOHdisJEhUSGllZg/jTf4/7nP51UGOJgpvK8zNxdYcM6ZWzum
j9c+w/acJX5pH1gLQmcoROYhBlu9pCdYUsevmQI9IpoQmYHHa+yWtj22TJbfB8U6
fgtb8oEjHFmNRp3xUCzcHwx3Q1CuK9AKpg3HXwGR0rbhhVeONy4pCE7j/IOVpGbn
DR4xhRRtkntnZldPdCb6FEh10XNQzGrev5H5SWrEm5K7e8iC9AoyFo299WBoyjrN
YDWbZKxA7ZlBEDkc7cZqmqKZeCgJGE2SKDA5ZYEBmWByQp5wM2Kuz9Z7xoJD3DPh
Dgb3bPgOBPyzpRhqqe8jHHPbh0orK6RaLY/9A3mD+r5clUh1p0RgsmrjwOgbJt6f
elqNTBf44BEQfHorBCufKXCiCSaQOHnMPbqWrqzKx9EDMaihT66AxbH61EIRnmQG
izjxvQyNN6XmfNDwbq5iQGmQYTruvgqJHzzjZzaNJyqNfEaKcBn2MzJqZjSp5G4l
18RLLgmfVy+CH3BABIrIbMBdmQo+3DAHy2RDin2SXDCEV1BC1aR2VNvDLicbKUnF
fk/oJT4G99ZfeChA6M95Uh7yet+iYkOu8mEaLvN0KtjMxYv0RdqMNXtWhvrPcScF
lE8b/riKa444URCf5517nTpJlNw8W+AKfkh3r0lWYNeC843hTMYQJJoKc8jUqguG
vYnbyiFSqc2sTm4IKyI9FGqOzryEQ3iJgdQUkDpnKtU+/KP23f5lQdY3eAQZpXIc
F2485ZwsZ15dUkfOV0Gh4l4IMZ3ulqO2n/DHgiQ8EfYvoLQVzNYc8CV5TjoAyAhy
BENRh+mTFKK8iyj8zTLIZAXD4YdKClXm7DoioXBT5psS5q2wrUjGSdQGybr8T2Uy
jP/znqAhW8stO2viNFSNFp/Bp8DN5/m5PyuQC5KtBNiF208mrtY3JRVWqI2KkPDb
ExZ826uAOwL2aq/vZ5STwZgrQdzCTAXpE8uceyoa5urGoTj+sv2Pdng8I/8pGkp3
3g+CQIXKXNvxPdG1xSGYCK3dOa9sxbl9Dc413SGlWiriaWCRIGIaJeptBXXlSb87
1fvgUHNDCiBthKiFk4nq42zNiDv+2RkE9MdQbpXFMyq4hWZCqu970cP8ivsUcy1s
0Bi9LWjbBU8L//BPSBsehmzojRnft86/5fyRU4A8BwU18hK3NZth29aaeUYyinxc
59OEwXSvprvHwWjehzOZ3uP+EuVnHg7n1QIyTcGsIJN82GtLSALbo/XUGvn8MuIN
tCZpTMJpfKLkYcWYqMZ6EnFBMxLq+q1sowSOK8luSoaYJEZ0D4JC7pddF5NbUWUa
GI7uFsYcSV4DoHVH6tmlXx16JwtOJ4eEtZ3rWsXtP39TRrTJs4/IdAcLVr9Dkfct
ChzZFmR8Yn0lHw6ybsdq+KIppr5RuEu2ukJUBnSzbJv+Ah2hnqLvpI4Dc6CZUDc4
wA+UOs/BXur4GQIG6DdlhdcThGfxV5Dc2uBuiDi+gB0/FGBE9AyTpHMz6jIPwi9l
B2b2z0EeQ3mC+YylTMW39eJTMs9FENPo1YwBBFBefrmZ7zkXncDI3gMuU5dYeDcY
MALpCp4S1Rd6bgaWh+TcyQiaAT4qKWXreAwyyQ2aaz6pfqhgZJcEsEOkWlXLNso6
pJvJj4rsaX3rOTTjOkxJwXXd3Kh2KfBRzFIllXBWvNOtPz/KWIQ+7MbL58dajAzJ
LoVNLOYtsVwD9BwwwoglkplnD1LYZAQvfORhRXyfLRx/ESjVqEcy00zWqMJe0CW/
0meTtoBAE2m2gSV5qK6vrH1WFV7OmK8At6+7fCk3Ifggn+Doobxzgwy5JKDO619p
sY9JMmDz1H8bVGyXSnjwccYkQynJgzZjBahhUIuINkcWhZ0wx19M0tlLkkj8IXlt
7LHnHRntdFSC+FhMwdBAJGoIHgHh+8iNZxis9rfOmHxc3IiJKF2AQihrRTiFd3nK
9OJSMdsthz0Sz2j1EPLrSCP26kadUV0ouuglzmdShJaXUNO4EHqAiSnSWEkN6kAW
+VoY9HEUIVXOZpVGes3NepxwcdZ9tDL9X5Myw6wKy8aj1qdE/Lih/lUWJFd41ihB
XpMfUgvaUkMhcUmIRYym8h9wMJ1wzHIX4jlXs2OoqrRd6DvJz67j1U2xZXOlrwXU
GkcZWNlY+oauceolOhoiJKsJc8j9fSKlSndjxHLGI7c16VKCo+551chFUNsOAkAQ
Qr0RWs19lHFUQX3E4XDhicj1nEDZKNRRQYXxzZnm9GgQba0s09J0xe9LgxB+YV+2
ts8r4sFkDRUOEj193/hVRgqbGYGOyE9e6o7qBOQGtIeMh38S2PU2qaMfzEw+GSGt
FJRyeuEIaA9R+66fMTxvVxKfHGim+dKDoSrnT5rWXSGpWa3eMP7X9yYer5dtqeD/
mDyLx0t/dryet/tf9Rk0/F+hTh4sDkfVZPJYqcn9Bz6EvfZJrdN+7IddUuAhg+bI
C9o0N1X7e2ZxGiUe55VFdnf04BgSuHm9upeWWAl4XnAOTMxy8s/9LZvQKR24Vnde
x+yN3Rmiftomsjg2a2PHxI0Ycv0LmgA5raQch9FshdNuJqORCWC1B86iWsqEXN5C
oUoUvpMMe0+D7+7HOQzG3fxsM1/mfLykCm0CWmreAVq5PVV36sdCd3gkj0unQfOn
b65BDKI3lAM7xNoEP45m7MesSfKMpel7b44krVgJg/IJXxW9N0xvIGe6biKUSDaP
SlY9By5znshYx4b+WVbG6dGFX+0dQf6AgBby1QbFsLtBQkJKm1k2pizAdT6fBKOL
YgbJlOom8MwIhvG6F/Vec06khxP3Yil2xYdxc4ivFso3cjT3IyZPxD8y5VQdR5HA
sdGOdJDyXjHNezvioZYGDSjwkFU3rXIgtiLenbaLz1/DWpbEZghxMM/gg/yfwmPt
U+nVv7kYyV9m9ZpiPTD97tD8Dfi1OxUs+yZq3FOS+bpqolyVuurvZUwbTLUpdfUi
Rdx9Qe9D4SdXtcGUVDfCdsWjTuvObIMd2bvC9ko6irEUp9eigGBB7/pXVKpnZq+9
wvbhXHEIHOwpq/HqWhama5nvaaXzXfw4HlvrNerzHUZLLMnCuahTLffgUN24c4Yz
t2cegCE6wbnI2PU/CQG1BR/JZyWFTZk9ZOUXPI4hiTmg/x8MsOoEtDrc0MLGktnF
t1oGOZkG1PkIo+REV00Pk47QfK1khspBo6UjYgwsBIbIHITKSOTQDF0oYEd7M86v
mN2swpYraAssttBCkAyGnYShxETX3a74nuRahzz1sjYjXmfLFHFOviSmLclyDeXN
V9XsnvTQHDeWbvJgwAEC+5vUGk6yOwB7T6zPh27fR3RDb/qJxpJPslPV/nNq4SR5
M/CzwD68rr2vjYW+eNvIJE9pUKY+iPME4g8qJhAyrSNUwwVsWWW9ue8v/t5EKV0i
BWJ8D6+sw3mHUdckT0SWQjzE7gWUz89UBGwt018P64J0gJTcy+Bj1JzrFvV59/Rt
C37ii2TmvYJ+Sd/7sfCbPQUKQFLRsnur0VjybsQagSLjNICxPN0/9qFmnGSTXtWm
WN0g6ZqdvYxBvYk9tDDTsOtrSHSPqIodwzJhov1cn5Sp/RF4p2e5UZKaOYsGaioq
lk7S6irCPemrrpVPZEUXJqt6atviTOamd4O0OLZrlYWXYQLEHUKNpjWifwP1q8eo
WNZiUITFLRmlv97/LolyYusXXGIxvinGG5JCRduO3rPSW9dvZrkBlsPhGH1q53Eb
zFlszZq0sG9Tb7Ic1qLioG0wgismN/6mqHuIjKyYwgQWNEG+jg1yvXg+S40GFudt
6mjcsEVl9hDmZC9G9BBZLbdV46lohCmwA8NkmjnvMIGJW10n3Wb9gJFEoMRh8SHP
ptKCOId1gw9Oy7RKrUR+tzbfc7Jv02QyYR+Zd1V7Bdt++16JNobyYG5SLFbm7F6d
0AxoxC5Dx6irPmXJpiYo7/WdiQbZubVVJiAp8c1YNjkwIpUV8LYZmE8cgF0Err4q
gNFF+Mrd62p+O1KDzMwjFMJ1Qz7v8rBWgm6vVg0EINs3eH0/k+Bso46AUwJLPXhw
aIuf/65qz1YcdpusiCfz1fbro3y2c41DbiKXMT3Afmj7n7Sw1wO+fy/t2T9og8iq
L4EabjHTgpg+w6HySWsiT0V0mfAeg2vZcZCNH4G32ZO/3neussJ3+agUlmXK+Zkk
5UTf43St+MalsnyGjbZ06ZDNCcWZyO4qDSy2MNydZHXu+0C2V28yTwBQ6b6BYeDq
zgQcqbV9lDtPQSGzIBLdzLEBNuWNDRPl++Ep9n1kbY4ZVkrtx+4JKt18Yx65s39c
cI6p86F/kuL77aX6W4GxCppUKmHpTRvfdMjd1rrULBG2i2x5oKBRG3IV5vsLMZKT
FJenUsIPCI3PzA6Z+X8HXa90zursEMjXCcvQuJqOciumala31SMwJzIKu5XXxFsL
EvQGcbOS6lqjOsjuOb1u9ZQu82zKuDRLiclo4yfKxAaXdKoFzx3h/Z4sE1TN1WkW
4opzc0oe2YjmNFYwRJf56YOGPGWoGddFu5gE6fLMhXnqJY03SqiFIL/kt4KnrTAo
HxadYI/S3ygLX4vcArnqQwPtsVM/UT6/AtwAZlXDJqVBGq0iSav9BF7MSsK2vQqL
GtdoBhInmYtSAvrQSSmHoaagckhO6v8DMhgIt/5R63UkFj+wYMsxe0zDhn/emA5T
F7gx10/fOSoYJPlfEwv/bQsB9BnRSBbZkPcADTt9u4hu06ZKipa1MlXXe8JJ4Qvb
k52QKVInXEvQyKTEPPksjjs0HzgkvxfdHqd9JNbNpUiIEaCoyO1SaNCb3tTAkv5t
imzyH3BGcmtXVPOfyJi71nckFjeqexSfcW0zoa/HD5QhJ11idhWtSAPOl1LPK6px
ie9NXJVdgOAYgbWvaXnRaQ9em/T5Kz0X61P1wajLUjFPg5BBDXXIT9mmTpEgVzaJ
KfLzGxs46U9TL7fXJJLZJ7Ml8ClfPsavS+8xAtQv7kctqCkRXaXhQpAkGNVSCdyf
ytfaWUSLkXo4cmeQDjPpsFYw9NABocIjPFS89V+3tHQYCyX78LsqItSJ9oQ5NL0a
gVT+YMWDc9FIGHWbCJCWaTQfSAzlTmOE9v0Kh5RP1A7YeEbtoK2CbsfX6spizQ7j
4DhM/Y4mrocfL5JXqFhNnIXBWzE2PM1ADd8JOHnqBqJNd8XeopZOfND6HB0gzKp+
HYQs/H4D0mCOyWkhplajp3yuLBBT/KQyjwVICXY7w1YyILvPPpeMVUm1WhKVKoAx
SsgCRHioMaczhaVTmxggZXWT4Ij0Ol09hAg6ZhE9w8nV7yp4Wv2xptNQgOgA55PL
FFlnNJEqdAT3FLeITZSNqVsJTQFwAXEkTN2wmTet1srG96t6DLobFjZQ4bieLFv4
YU6YDf/fxMEOGNdQTY8ed6WB+hkM2kceBSbtWes4CFIPMxz3qbkw6zkPSG07tv94
dm5zszLJT0ogFcHw3VELxYF3nCbK8F9hy6fk1m92JDeUWVNGDJdo12NtKupht2/W
OC6TVPRy1aFM4gZS3A2ng4kzuMsTevsH0fN87d2RfeqwjwYgQewxFfkFouJw13Pu
XAAEV7GPupmNbut99UTQqEsoaZCUUC6eHfHVyDhzzdhBJ9JlgZ9hxXyfIEROQCpk
P4ed8iYE504ePN9LKQUU+QsnsyvQBYQTlJut2NG/BfWfLAvVHWhFZbqaIGLGgz8N
4aim+purEpoqrSw9jtb0g1qFGMgMIUiRx8mm4lk7MoGVmbzdXY6NvKgtNV7FTxsA
lHSfNjiNrHjvVQp9NnVnio724ciXe127dICuQ39+Nn1oSgM5YL0PS7xp+Sc94C90
60X6wAqlEy0o+7o9cJMUOpdDfjpA/eMExVZwkV96nHF5jkNctT6i4J0J/v2G2Mkz
cAhbWGJkzMc0uSVvPyx755u44OlOoeBGSmfwh/CrR88q1zkiDLsWqF5SOTvruGDj
qKrTd6TozJMHnD1iJvjeKV+6S70JSgYXmeJae5IM7HHziPa7N1cY/Gker64HyFqD
deu4E0fQ7g9/wfxpFKh1DjDMFDYriwb70Zp4keUoNFEhGu2en3uD4bC7aq3onjIA
3GLdnE6KLpHeNVqODExwqtEaD2q6+J5NMQzn83k/Jsh1/Iy8xtPKc4SqnOqfDvLZ
kGCxIwGNdHz9bZhJfaCGfuAa1CZjKkuVbYT4v8dzfVi6av/ii/5SOXU5Tklb926u
DhjCIVpzRHwpkTNMAjlQtrJFA/SK7T6faM7suP1tYG9lphRXZn7XF93hDvZWBjUU
C8xQePDx5ba+y6NAui6gTXrySw80YszsgRKQYCXMyOtC1aC2IocWtPcDK7QmvVka
DQXFW4Ne7Kau5Mm7QQ9wIic3qu5ZWBSMenf7Aj2zbfiOS4V/3F23KgvSd97yzCaD
5XuG2paYVCzA1CpJbRxU2NLJ1keJ2jP20BDhc1OAFJSvlmzClJ0RSyKZ7PKH6384
8JY+KwUrYkmqe9A8A/chl+rRgN9JSalKYuiinkyN1h1ZNmmsRqWpFFF6AkwMYlBA
2YFYThZrpc2aHhsXL6ezFsTZVsWmLPWidHboeY8UJsUwNUWl/lOnaggJ+gP+fkOY
jm8Z4SDMEqNGRkYvrAA8gTlNz1CLYk7IVpHNo58IR3gQSqij9/kqCRKaccFUZ4Xq
kSz40sBzwIsl9cacznRdD+5CTXVVOwKwkVySIoVF1GlQmVl4wHj8RXBHnbahrS3N
DywPy9eViX9HG4o4oUBscEnDgQjkjRVbMxS5NLPH5SLy+8I8+WCZDxiQTbE9+QUb
x08QHZgU2BJBLpzm798lInqTaLSUlA5661Pv3r+X6ZgrJa/R5fjLLi0Cseb7mlyh
gEPGnS6fHCeZSlU6B4cz2CxE3XeBNUTjrN9uYN5ilGJ6bv88at0q2hykSrCe2mJ3
aGovcC8wPCzM+eLnA0MM7oDQKrKgRKO/ZVaO7mXrYrFIUVhh4O8ddl2Zaa0QGIhF
OloaYQDlonPdrdZjpr7nhjhr+HzLk3mdSr1Ge93TXglcP0TwZrIs3Y3yN5TuvO4k
mLL2wT82DDv85ofPBxQ75aPFsXNlq68sFHkQ1VgnspTpDLIQO4N4oqyPKVizUOsX
Zh9RGgWra+YvpVYmrqRZkGyricBS9tgKIjRnST/7JuWBAPB9BnHg8OsxuyBSMfSc
3liFQCISw7AgW0NZa4Af1aXHY5gHASTuL1qEF3XmO6R1S1ebp3dHEMEpqW0BZ8pz
Z6OOeRLPjE/IfOXEKaeU/AqSBiaWHSDgVgyW8fIVO0nrHDUGA0WPgxG2fpN/zqlc
gIB6ckTf8jnmz3XNxJa190twA970xdUA6KhIzHvQSZnHAvyI9m+OOMwq9WzNI5aH
cVIzs2503/LZGAC3qeiKPdaXLjc6SuMRuSIHbjeZfF/1+4GPeYnyKg2sWvqUFpzQ
2xECbuUzXfjzN7USGxsIWRbhfrbGqS0SN9XW1lvDUSqU7hhyv8qdEMdO/MGYFQPF
ZGzBeHbBFZdb7Pmp9mKBtlnbqRTZKracSnZN5fWvwtpC44ByyAWcx8NSWGaT1SkR
Dz/Cg/+w71bl5NpJimDWcoWVwnNsxLrPWt1M9P/+NumzjSOPbsaPhI3eG2JIowAI
vEv0+e1esMJcL8lqSWmw/bhRhmkT38iNCwsb3tywm7kfGouXYLeOKl88PWqLq4Ph
x0JttTA4gsjodxzMsa91HimxD/FXVEKhmyWu/rFYqaYLivrblqn9is8wAHx2b1dU
kW/5/NvPKs2AgfwYQT2bFKQs054ABSP9GJ3erXDs0ArNpzKdmhqThgoRYXivg+Qi
ifxLLOGNr55qH19WxTOvt4eHI7lnpY1IwaFoz7mGjsPmfsmAPAvz1geKRdlzXZdX
VdHCupKJzImC8L/2A/b8fopfZuAltEDgxzcATDrKQjdIwShX8qnoUnLkFWRmYNKm
23d6ZyvKVtVzszgICppGjas6Zaj/FalZiXSA6zRVmfzSMlTpG9Rw4WekZyZ6ySyT
BbAaSUqdfYC8aEb+sNDY/molTdSt7MAU7YiHoY8IMqchT9KocYjSvPJHlBa4bAUE
4mrBzeFC+4oWw0fjPyGHFOJniRSOLu7NJUXJpsuA6HfN7RYCGOtIzAf8MK/QVYeo
ggDxN4MC/SMhVBdjtemv6IQaflJce2MQaZwQxKQqQGayqNKB2T2wUg0ayr3ylFAy
bFSklJqTRVUj1lw8X6TcvFLOtnt0nXW7T32OLYkFz/H6IpAaGaWvuMGTTC2JFOtQ
qf/5f8iJ2lJphEj2gopZQ0yCKu2pjBmbTdz8f9EpKgsEHPM49eMuxa1jgwomOEfz
XIdrtB2AFAwrxGkGj+/UD/A/ezzvoDkOmKXOIoizU4vXInlM8niy/Sohl5IJ/rwm
nvLegX4wgjhA6iVqlXJ4blwokJO2CACMmtBywjLkNmttXt7MX6uFhECqRm0AVh4C
O9gvK8E/V/zFQt9gBWw8urmihyV134fJx+6H/z7KnyqqjhZVshWY40xJcriM3Ir5
Km0tUj51sjrfqPb/RagwDpU+P6NouDj4CMc5Y+OrnYowZm5kUNrguMmFN9Jphk9z
wYqzl0rbBxi89P9kP2IHx864Dj14ieE1Fdw0skXru0XyuZf29JGPBRdta29XERdz
kampsu38dcBfqkxZEnTlQcg+x8XrXjFILcUwVZTVdI6+92oxuJ4uJdxDdSayDq7Y
D+dLKsTfKKRkVN8l0ekXb26fTOp3Hkr72TTpMZuIggAtIWEbDaFD0fpw6/yWsKU3
xMph7MeRuMPsB6GHZvqYMfB23PRTOrSzOUpDumozRhPoQY0hyYUFxlF58/PMajM5
VW0vbdb9J/4U9jTq/Gi6zFlqcS4T6MxNH/QjdrphtGQly1sNb3UNVaqLbTkQoJa+
UdeUyc0oMKwJxAy1+O05xL+pnYPB74Ozo5zXaANNYszdp1ZcyRaCNc4PuNbmZzwD
hYUibRLtuYlFPnn28wY7qaqbUUjZ3qi2yXXaLeHJho/1TCO0omZMSOYdFq3LdQsb
nLsps+BkkfOOshnz84CZopTrR4h5BN+6U/wh3HxKHRhobXuJVjrz6UM0qEayAieI
/t8T6pOhKVz5sxrDkV98wGyke0z4DEl9eN5HWMFruDlCe10Q/I40QOM14Dyi7PXk
jghTcXTiAxMAK4UeInQ6v5qFTpMd1BvrB0sIwXc5nAb7brXzL+MqQIsdOfrgUinL
4dnDA4RKk0Jrzeki28+PzL/1MHrT1l3FehBzVQhL9xmiJPXe/DfMvy+MVjPrZEzy
rFxNvAyUe1RrubjgUMMwJKVrGdgUW383XsjUr0kZ/SxI5ZTH+vfDJTSUeeBByBA1
eHWcBAMvmAFMj5B86+ICs7yBqsWmoln2GgfYSOdDKSsyYyB4kqFLKrNoRJx19OfZ
KCjNdfeNrdhEAOFYoyunE0pY3s+Ev8ga9u/enCu5coGU1peLW7U6JA+dXTJpm93S
PxiHkw7ss9Xqey6WbWTDFyijkdnE3rA8CWxlTQ2zpiKbHmbQVNACqfYaXxJgqFY1
luvawURUW5PBKOeCuuMj2/tDIQoxtCQwi97N3dK+KuCD+tZ1QiDSreSbVTZc9Dke
AZ1EXkNFgugT7FkqiaTBsYbrdJyRsOujQ6rjXv+t5Zfev+XJUCB0HW53Oj0WLndF
TOY6zWjGREfYTmC/Z1y/8xclsEx6ZIOqbUHsYej/MVK3hG4IzmXLf1a2vgQQ/f7w
FltE1ATW2w6devUm/DzKkLhhlk3SXCcARpobtfkYVqjoqKUqLM21+vU/M+Dd49QB
wfMjx9ehEwwy5lImozrSE42Wl4eFdMfaC4296dQtkb51sgkyVlGN620eNBSP2sVO
xGIyaNDF0/NZKMcxLv77ML4y7bw2RqA3thtQjKEdkXdDvp285vrfvroZSFoqU9hF
Pt9mUbuBkbEl9pF2Hb/f6Bcjk+HLBEPNj5exH6JaR2+k1Ayd/UBKP0efkkw9h2RL
RMc+KwqvMSYqX9YqjrPKk6flXoRiFibHc8x4xiJuwmJxj9B5rqSfG2B4GjkeSsLy
pQj7Dbjsp/iHWZ1FhZrXrkrOkqm7/zp7PazpmTewvOYpmoRdWgKD9cuRHBI65uqE
K5jjFSpwrv+26+q6tlJJ4wbn/6dFS0PE16SKIMI7WmYNFy71ZIOV6bEHpzT/0s79
9jZLG0XQ4fHcdpvsAA3nD8wK+OaiA6acIIXASWSQx163EbulDyLl2OmWAz8xV7uL
yy/TWjO2s1YFLVJVwzGeqFUmPtjO0PP0l/94Oe3a3NkAxOnYl7Che3IDuo/cZr+y
Z99txTCSoaKpetSKemWFZIjrmqKBWU3heWngzJjrSGi+vVFbMjeHED3ffXfl4pAA
`pragma protect end_protected

endmodule
